//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.10.03 (64-bit)
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Wed Nov 27 20:13:50 2024

module GSrom_test (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [14:0] ad;

wire lut_f_0;
wire lut_f_1;
wire [30:0] prom_inst_0_dout_w;
wire [0:0] prom_inst_0_dout;
wire [30:0] prom_inst_1_dout_w;
wire [0:0] prom_inst_1_dout;
wire [30:0] prom_inst_2_dout_w;
wire [1:1] prom_inst_2_dout;
wire [30:0] prom_inst_3_dout_w;
wire [1:1] prom_inst_3_dout;
wire [30:0] prom_inst_4_dout_w;
wire [2:2] prom_inst_4_dout;
wire [30:0] prom_inst_5_dout_w;
wire [2:2] prom_inst_5_dout;
wire [30:0] prom_inst_6_dout_w;
wire [3:3] prom_inst_6_dout;
wire [30:0] prom_inst_7_dout_w;
wire [3:3] prom_inst_7_dout;
wire [30:0] prom_inst_8_dout_w;
wire [4:4] prom_inst_8_dout;
wire [30:0] prom_inst_9_dout_w;
wire [4:4] prom_inst_9_dout;
wire [30:0] prom_inst_10_dout_w;
wire [5:5] prom_inst_10_dout;
wire [30:0] prom_inst_11_dout_w;
wire [5:5] prom_inst_11_dout;
wire [30:0] prom_inst_12_dout_w;
wire [6:6] prom_inst_12_dout;
wire [30:0] prom_inst_13_dout_w;
wire [6:6] prom_inst_13_dout;
wire [30:0] prom_inst_14_dout_w;
wire [7:7] prom_inst_14_dout;
wire [30:0] prom_inst_15_dout_w;
wire [7:7] prom_inst_15_dout;
wire dff_q_0;

LUT2 lut_inst_0 (
  .F(lut_f_0),
  .I0(ce),
  .I1(ad[14])
);
defparam lut_inst_0.INIT = 4'h2;
LUT2 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(ad[14])
);
defparam lut_inst_1.INIT = 4'h8;
pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],prom_inst_0_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000017767;
defparam prom_inst_0.INIT_RAM_01 = 256'h000000000000000000000000052492B2242492B6C8909248DB2242492A6C8909;
defparam prom_inst_0.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_20 = 256'hC52A46F806C4D98788C75D9FBBC21D2044697BD0F17CC4AD4DD1D9869675FFDE;
defparam prom_inst_0.INIT_RAM_21 = 256'h578EDFA38DBE7B0FD33589F7FB305E28DC712113DAA265CDD3A6E50B98265ED3;
defparam prom_inst_0.INIT_RAM_22 = 256'h898F9DC65427B02B7D0792437D5959BCC9D58E49F430A561F101CB3CD2B3C39E;
defparam prom_inst_0.INIT_RAM_23 = 256'hE0D519075C8CF5F0AA8BE6301D01CE2EA5593BCB589A34801435160A3CFAD69D;
defparam prom_inst_0.INIT_RAM_24 = 256'h7ACC9A99FA79159E696414D5330AE4BDDB8F14F559AB5119D43BE19A22F2EA89;
defparam prom_inst_0.INIT_RAM_25 = 256'h380F8CA8B22D0C07B3C7783112EF57211EFE8B65C9D0BAD72C5D0AEB32575B85;
defparam prom_inst_0.INIT_RAM_26 = 256'h9B28C4F697A8EC6950020137CB796057E41F9844DEB0CD148C992DA249563F1C;
defparam prom_inst_0.INIT_RAM_27 = 256'h799494037054607B1C29C8BF9978B4B3BFD571059297500439F73376B46A504D;
defparam prom_inst_0.INIT_RAM_28 = 256'h11C331E95E7C491DCC9E19BA5B07F3E7A908F28E8EB1979D0ABC30010880B506;
defparam prom_inst_0.INIT_RAM_29 = 256'hEAE2A9C403F6F259EED2AC6EC28AF7D16DB6B4A50C130C87E3B9B3A05342EE5A;
defparam prom_inst_0.INIT_RAM_2A = 256'h40578B79D0C6E0EF0B02FD27AA541353DE43CEDF24ACF0D68CEB43719986454B;
defparam prom_inst_0.INIT_RAM_2B = 256'h1939DB4A6D233E7294777025B010380364975591C1FAD29F6FFA2BF527719899;
defparam prom_inst_0.INIT_RAM_2C = 256'h4127EB3311FF07F7593FA3F9576CEA70A142B09FA37AC8D118983E84B8E5DCA2;
defparam prom_inst_0.INIT_RAM_2D = 256'h9A24CC37BF7841DA0F04F4A5217CB5C078B399EDCC4B51382838C2FD4F20FDE7;
defparam prom_inst_0.INIT_RAM_2E = 256'hF09393D8695AC9A30B8E64D8C85BE120D600F4B553E3D74AE61638C5CC56A97C;
defparam prom_inst_0.INIT_RAM_2F = 256'hBCFE7BA4814CEDBC148AB46966ECB0CEA2A8B5F96DD10D1462CD0324047BC236;
defparam prom_inst_0.INIT_RAM_30 = 256'h96A87F9424796DB105787EEECDC706BBC98435CC25424981A8D6595B5598B56D;
defparam prom_inst_0.INIT_RAM_31 = 256'hE2F7F5B9D2F7CCB71FDE134199048299CF7C4E7E687199559268003CA58244E8;
defparam prom_inst_0.INIT_RAM_32 = 256'hBAE93903E7078FDB6D64E780502073C31D09BF782CC2F0417B95E5F8A5166B24;
defparam prom_inst_0.INIT_RAM_33 = 256'hC3F8AFF640605D2C001FEAB0F50207691C58E80331174101FCAF1E59DF51EC83;
defparam prom_inst_0.INIT_RAM_34 = 256'hA2B4D07E953469749E33265FE546BD12ED5164D4015F20F1BB5F0447F94FAA41;
defparam prom_inst_0.INIT_RAM_35 = 256'hF62AD5D8A1AE0B155CDC42C8266F5C69BE2C7E2438BC33D4D21869D13F5B95B6;
defparam prom_inst_0.INIT_RAM_36 = 256'h89B2E9166B1EDC484F90A0E5F503BA1BE4887A59F24723EF412531C02CEC5062;
defparam prom_inst_0.INIT_RAM_37 = 256'hA5E64EC4F86E514A609A156DBFFF2ED4E09BBB591969FC8192AD7F3311E22BE8;
defparam prom_inst_0.INIT_RAM_38 = 256'hD969291439A738A16D4EFDD7961B1F4539A88EDBBC734AAA83B8A445F923FDA2;
defparam prom_inst_0.INIT_RAM_39 = 256'h99F726E9955C337A8977DCB57EA31ED7373A9EE0B20ADFF75D5CC9DC51B0B3A2;
defparam prom_inst_0.INIT_RAM_3A = 256'h818A405DA9B4F1F97767EACD397F1E69437DB107247266B858F9A1F435C39E0A;
defparam prom_inst_0.INIT_RAM_3B = 256'h99003CDB61730B190AD1B4F9E5F69C52CCB3ACF0F136C06C36CD311FCA208BEB;
defparam prom_inst_0.INIT_RAM_3C = 256'h0BEFBEAF19DB0ABB7F6D35E7B63DF2CAD991096E48BF5F5499CB439DECFE67D2;
defparam prom_inst_0.INIT_RAM_3D = 256'hFB3124BF940A5EB3D9E3C28744A096C15F227652DCDFAE58B4414CD2289AA462;
defparam prom_inst_0.INIT_RAM_3E = 256'h99EBE15634E3E8FEFAB36059F9D1CACFD3D3ED6504ED2CF277C095BE857494CE;
defparam prom_inst_0.INIT_RAM_3F = 256'hEB3C43BC2882520DEF036C190B8FF6DA45FA5D7B7D0E7FABEC279950C2286830;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[30:0],prom_inst_1_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 1;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h5E0E932D62557ACF857FAF2E94F3E942155BA2B5DF23F0A1E270BE41215AA4C2;
defparam prom_inst_1.INIT_RAM_01 = 256'hD9CA20E558AC7A19BBB49F4FE27DC1894CA86BE9A51C82BA66D5A1C506DEDD3B;
defparam prom_inst_1.INIT_RAM_02 = 256'h00CBA6F76B2179FBD9E6FD4717E3B9AA58858EED79EE101977B454168A624445;
defparam prom_inst_1.INIT_RAM_03 = 256'h2C237B2EA161960D053ACC043A5BDA4DCD8B17719EBE48568B3A94FC3FE8D41B;
defparam prom_inst_1.INIT_RAM_04 = 256'h3EF151535E5F5E1C2ABA902051DE0F62303AA37BDC29757B70C9CC7094EA7AA0;
defparam prom_inst_1.INIT_RAM_05 = 256'hF283A5C4DBFE0C343F222796C9EC47A788848F13BEE6612E419F0B1170095363;
defparam prom_inst_1.INIT_RAM_06 = 256'hE7532FFEDC18521462288E7ACB65E1BDD15962617B505B85009001150B931BE3;
defparam prom_inst_1.INIT_RAM_07 = 256'h6C744CCCFD17E49C26681BA1E69EE53D330B8533D57161E1DD3465F6CAE4B0E2;
defparam prom_inst_1.INIT_RAM_08 = 256'hE8BE3018AC472C71830E94A9963E05C5AFFEC967C76A9ED9995448850BDE9245;
defparam prom_inst_1.INIT_RAM_09 = 256'h61CD683BDA410012B8009CB5C1E81FEF80BC1685C007DC7479F407839F6C39C1;
defparam prom_inst_1.INIT_RAM_0A = 256'h98C2B5406C265BA4241E4E5B0316DB1E043BF80CA42313655D72995230DDBB3B;
defparam prom_inst_1.INIT_RAM_0B = 256'h4FB4823127863426D34A027BEC3BBCCFFB7639ACFDBB841C29C8A5E23F50A2EA;
defparam prom_inst_1.INIT_RAM_0C = 256'h9FF38783AA2FE5DC68967DFD26F07F30F17CD47AA0F99DFF2E0B623519F8B329;
defparam prom_inst_1.INIT_RAM_0D = 256'hE544B73C3D67911174A2F144BF8BB7FE908771FE5C30913E3D79C8D9D5406102;
defparam prom_inst_1.INIT_RAM_0E = 256'h2871F66DAA6792A07942C518E4AA8484B34654B1288F5D8B440CE129DD9C399D;
defparam prom_inst_1.INIT_RAM_0F = 256'hCE26F7B9E372CB701A62E21252B9C4F1419DF58E8527F7BC64DABDAE167D70E9;
defparam prom_inst_1.INIT_RAM_10 = 256'h9165FA57E0A305107E4EC68C45BDB916C83C672FC8BD60E95024F7D9A5751624;
defparam prom_inst_1.INIT_RAM_11 = 256'hA5E451A3A7611098219F0FE8D3A222F5D2883164DE4F686007EE028811E20655;
defparam prom_inst_1.INIT_RAM_12 = 256'hB9B5CAE05FC077687473B1AFE7D320B7BC9AAE3E23ABF76AC484BEC2C76E491F;
defparam prom_inst_1.INIT_RAM_13 = 256'h15706D8C053CDE2674C4270562DC85DA6EB422B429BA18EF7458E6F390712806;
defparam prom_inst_1.INIT_RAM_14 = 256'h3DF5771EF7785ADA16AA503121B419725764A60EE446A1A68ADEC7D70CEEBAD3;
defparam prom_inst_1.INIT_RAM_15 = 256'hDBECABCE38FFE793B925EFB4D2000C98761BE6410C12B4E6F466EE7804970CF7;
defparam prom_inst_1.INIT_RAM_16 = 256'hFC7980001A7F81B4674E98660FFFCDCA03F1CCE1544119DFE1FFA0BE7B0C8F2C;
defparam prom_inst_1.INIT_RAM_17 = 256'h85AD75A42A83B31F61FC7C15C4B305B49DCFADDAE2FE1920FB0A00101BF80550;
defparam prom_inst_1.INIT_RAM_18 = 256'h4DEE50D1F84F9ABFC9C628D0F102BEFBFA5F42204AC0EA0024B08D9B97801A6A;
defparam prom_inst_1.INIT_RAM_19 = 256'h415A8EE92F1ECF0948D727E079AB82798A45DCEB752EF11A18BADA75CDB7EBDB;
defparam prom_inst_1.INIT_RAM_1A = 256'h7D2EA20F36C27C58FAB8895CE6E6A87538DC887969096BAA5DD38FF5D4F752C1;
defparam prom_inst_1.INIT_RAM_1B = 256'hB445BF6C83ED712F346CBA65ED8CB0BB3F4C2607A5112E3EA76B924BD6C3A8C1;
defparam prom_inst_1.INIT_RAM_1C = 256'h2786FEA0E36771F38588019C7DA3A37B1D2C84695A03E556840564B5A5EEA81F;
defparam prom_inst_1.INIT_RAM_1D = 256'h21F4275F31CA20D14D081F90B16F80FF946343A2DFD913310CBFA2D5D7F07471;
defparam prom_inst_1.INIT_RAM_1E = 256'h4014014F8D90000050001E948007E36400108002000006DF069C3D317BFFFFE0;
defparam prom_inst_1.INIT_RAM_1F = 256'h644830218482000038A1C9200130020002A4E09810FB5F6C0000000965FDC800;
defparam prom_inst_1.INIT_RAM_20 = 256'h71139BDF3F2E900148FCB1FBD7289737932527AE8B32C202D410FD0000001020;
defparam prom_inst_1.INIT_RAM_21 = 256'h72D73F18BE3A49AD44D1FE051F6D6DBB3CF027BF146106FB3A3C450039C4E2DC;
defparam prom_inst_1.INIT_RAM_22 = 256'h33BD17B9D4548141A80A64B87B6B9FC1A532FD215B62DAB6AB383923756FFE2C;
defparam prom_inst_1.INIT_RAM_23 = 256'h070420B20870A19CA5EA6F576648A051D99F16B46BA80939A824472D86CC7B9B;
defparam prom_inst_1.INIT_RAM_24 = 256'h62542E24DDE77844A07CA40AD23991EF861CAD250117D1EA06B574091EF2DBEC;
defparam prom_inst_1.INIT_RAM_25 = 256'hDFB9AA6EAA5F4E6485E6CA4AAD1FF19F1635B357EA45E1CD42B51BE48F3A3765;
defparam prom_inst_1.INIT_RAM_26 = 256'h4FD1E3D168CC202D2E1E27707E6B840A315705350DF18DC9A4BA58F3783D2495;
defparam prom_inst_1.INIT_RAM_27 = 256'h0AF1A9257E3C839FEFE6FDD00DD1BD6A7D8617C0A246B2C4B8F50C3B36F7B05E;
defparam prom_inst_1.INIT_RAM_28 = 256'hB536BC7A48EF7497EB181FC1E095A89CC04A4D797F749CCDD2F4008E53D4A40E;
defparam prom_inst_1.INIT_RAM_29 = 256'h31769CA8028154A8C5C21DCBAF15CA09975E127F6FCA9155C0DDA891C7FFDEF8;
defparam prom_inst_1.INIT_RAM_2A = 256'h19E39919C34240469DB63AA6FD05E84789BFDD1E476239B94A738624BC0D78A3;
defparam prom_inst_1.INIT_RAM_2B = 256'h6B5F0B13D5247F2105B9EB532EC4D080CD679E45E04F56930A289AB0EEC7FFCF;
defparam prom_inst_1.INIT_RAM_2C = 256'h7FF21F673FEFFF51950CC69649392C6945461931935C15D7A318AFB7572272F8;
defparam prom_inst_1.INIT_RAM_2D = 256'hA5475F14E8A8C213922F4FE667F56D0F6EA339D23736A99F3B389E0D29863891;
defparam prom_inst_1.INIT_RAM_2E = 256'h102D2B3D68802DA79E75786C6B822513529D68EEB022DB88AEE5F835C341866E;
defparam prom_inst_1.INIT_RAM_2F = 256'h174B7179EC73FA4FF02D4D1308018849E87B36A5478A18CDBF167A6F14310E32;
defparam prom_inst_1.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000001E79E10;
defparam prom_inst_1.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_1.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[30:0],prom_inst_2_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 1;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h00000000000000000000000000000000000000000000000000000000000057F7;
defparam prom_inst_2.INIT_RAM_01 = 256'h0000000000000000000000000186DB39CF86DB91E77E1B6E039CF86DB01E77C0;
defparam prom_inst_2.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_20 = 256'hD37D41C9877515AE20FC01E8B27C4E2366DF1C85F1AB45490C2E10D4B457FFC0;
defparam prom_inst_2.INIT_RAM_21 = 256'h4AE3E083D7235F39F857DB39A79196CE8D510B0622304B0A6C7BF7D7EEF83BB9;
defparam prom_inst_2.INIT_RAM_22 = 256'h6662C3C2CEE3A319A78945A9801314A2BA58016549A5BC686CBA7177BC01878A;
defparam prom_inst_2.INIT_RAM_23 = 256'h26D187A7BBB2CAD87CD1F0476D1C5CA283733C308A23E09115D8065D58F68DD8;
defparam prom_inst_2.INIT_RAM_24 = 256'h6E59F647861B3380572FF230F1265279BFA0C26CC799536401BF5529C405FD20;
defparam prom_inst_2.INIT_RAM_25 = 256'hAD4F3C58719CFFF8DA97E60F0E233F01D45778E3C73678284AF606670E31387A;
defparam prom_inst_2.INIT_RAM_26 = 256'h78E83C1E7500F0926F9E06F0C706819A4806783C398FFA192918E3A1C731FFE1;
defparam prom_inst_2.INIT_RAM_27 = 256'h593AC0385ED5E9460CA2E857E3591184FF7AF0FFABE679FCF80DA0F1740B996E;
defparam prom_inst_2.INIT_RAM_28 = 256'h7348D4CD78A2EA49CA9B1FB9FFD746CB0A1D7B0549F91AF07D094F1C97F80A83;
defparam prom_inst_2.INIT_RAM_29 = 256'h596C27F2B2CB6B02AC06BEA58C5973E3D3784FF23A0E833BAA0A01479369CB7E;
defparam prom_inst_2.INIT_RAM_2A = 256'hED103B3165EC69DC6100E5A1432CD4BCC8F5F557C2E3D37224F64B85D2CEAAFA;
defparam prom_inst_2.INIT_RAM_2B = 256'hABE8328D5B25998479EB71A3BA54C4DE64B3FCB9290287F579CE11160EFD9B89;
defparam prom_inst_2.INIT_RAM_2C = 256'h713F25F40C849AF53C43BD9B14A995A351D907C1C3130BC1AF27D54CEEAD9CC2;
defparam prom_inst_2.INIT_RAM_2D = 256'hE29A963FFEEAEB28A87806664D7DB3A8951164540A0D9E3D66A36FE44F016D76;
defparam prom_inst_2.INIT_RAM_2E = 256'h0031E5BF4D9A2756A7FA7985F2C34A3FB2AA532C60E41AC34B91E452A41F3087;
defparam prom_inst_2.INIT_RAM_2F = 256'h6315F6A12B3089C38C586C749E8125BF34C0732B2C1B0C9275BE25C4732951C2;
defparam prom_inst_2.INIT_RAM_30 = 256'h7199E01A9584247E18781DDDBDEB6CFE9B8739FC1CD92014650CAB2399E78CDB;
defparam prom_inst_2.INIT_RAM_31 = 256'hFD0874787006693F33801C0078C39FE295832600707078CC7072AA7DEC7C78E8;
defparam prom_inst_2.INIT_RAM_32 = 256'h0116C6FFE0FF80207184E07FFFFFF03F03FE339FFC3FFFBFF8741FFF366018E4;
defparam prom_inst_2.INIT_RAM_33 = 256'h7C00AFFFFF9FFD03FFFFFD40FFFFF896FC07E8033E17FFFE0000FE07C0AC70FC;
defparam prom_inst_2.INIT_RAM_34 = 256'hC275011EDC9DC585804CF1249E5196F7A4CE871401001F01BBFFFFBFF80055BF;
defparam prom_inst_2.INIT_RAM_35 = 256'h1D199CADA1CFF73997EBE4D147B53EDB3B3750613B690F324E3B2BE8688C5844;
defparam prom_inst_2.INIT_RAM_36 = 256'h078E670072549C243010581CCCC32AB21DB80007F1CD6FCADBBC97C0037C3529;
defparam prom_inst_2.INIT_RAM_37 = 256'h6CDE003BF9D9DE6F2AE6C31C0000E9B3FCD11584B4E00080719C87A5A6E11800;
defparam prom_inst_2.INIT_RAM_38 = 256'h6AB11B73F9A0F8671F8B5767B278FF42F8647F12EABF26678007A1CC3E35553E;
defparam prom_inst_2.INIT_RAM_39 = 256'h85CEEB2274D3FB787D0E3C19B4330630F73E81E66DCC9558333C3FFC30738C3B;
defparam prom_inst_2.INIT_RAM_3A = 256'hE8AB307FE562EC1D9B785EE1B84EE9D9D37CAE33EFB4446530D070427EA8658F;
defparam prom_inst_2.INIT_RAM_3B = 256'h33417E6A2BDD39B87858D192850D72F6147ACCCBB704BB5907AB55EF5326E3CE;
defparam prom_inst_2.INIT_RAM_3C = 256'hF35AC15F27B6F838F809629850E34E71D981FE7522CA760C3840C77B437A7239;
defparam prom_inst_2.INIT_RAM_3D = 256'h00EB1BBC73E9CB3158672679C750DBD6616EF631C03FE06294E1C2311870A061;
defparam prom_inst_2.INIT_RAM_3E = 256'h64933ABE660AA4A9C450F2A23B0EE9DAC33CFB1505FED1A98D78760D87025A95;
defparam prom_inst_2.INIT_RAM_3F = 256'hF9318CE3448CB650A312A31E809A96AA24A60EEE66A8887B34B77FDFFDB21A6A;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[30:0],prom_inst_3_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 1;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'hED23B0FC2BAFEFE6BD149F44B1CD0E65B5A59225775C3F0922C535D6762C73B6;
defparam prom_inst_3.INIT_RAM_01 = 256'h9BFFC2E18A5AB839410F9328DD79A1F8BD9EF3C2F791FDDCB18109DA9F4CD2CA;
defparam prom_inst_3.INIT_RAM_02 = 256'h99892A781ECEDD61240FC29B6ACB072FDE21AB73D1C5A0F5BF9C0086E59F667E;
defparam prom_inst_3.INIT_RAM_03 = 256'h85B49E2D23CE0E128EA96D0354A644963D274EC2A1727C03B5FE6711E3C94CD2;
defparam prom_inst_3.INIT_RAM_04 = 256'h0C79DCB83C74E5E853CC89E2D3176BDF4451BE9F664621E5456EE063C7E412D2;
defparam prom_inst_3.INIT_RAM_05 = 256'h288FCD7BAB5E162D6253CD4B9CD16C376E73426CB5AF62AF2A9B187E71EDF0D8;
defparam prom_inst_3.INIT_RAM_06 = 256'h088936EEC854CC6627DB752B5C4AA7AA3452F44651717BF669E3D0A94F1F2461;
defparam prom_inst_3.INIT_RAM_07 = 256'h492825643E601DF81E21D9DCD215A6060D047C9799A4974B640E86EF4496597D;
defparam prom_inst_3.INIT_RAM_08 = 256'h0F383FF883FF2C0F9F0FE70E183E7C625003C748067314E7B4CC0E02F83FF246;
defparam prom_inst_3.INIT_RAM_09 = 256'h1E64D4E733FF001007FFFFEA01FFE0107FFC017FC007E07F8600007F8093F83E;
defparam prom_inst_3.INIT_RAM_0A = 256'h456F13FFF30A76B1B3B8FEC08D9E028F6A2497E575F82831E79A41FAAF543B6E;
defparam prom_inst_3.INIT_RAM_0B = 256'h4F3F0781A6C9F77D6A6EAAD0C0A582129006B01105940EE5BB94E0F486AC9884;
defparam prom_inst_3.INIT_RAM_0C = 256'hFCC4DCAD62586295E2054AEF04660229E9C80B566ADB7A7FA4A20E0A506637EA;
defparam prom_inst_3.INIT_RAM_0D = 256'h7507E87D2F4981E92A88B3A5B3C3441D318DB9856F018D2C7AA5052252275A6A;
defparam prom_inst_3.INIT_RAM_0E = 256'hBDFDF6A483229EA19A62813F506D3F309FF692838464746D521ACA2C85509F91;
defparam prom_inst_3.INIT_RAM_0F = 256'h17BC3C456A9095BBC0DEB5D16574525DB4F717C61A66AB28923CCBB2EE8D1512;
defparam prom_inst_3.INIT_RAM_10 = 256'h061C19D01F365A6DB3D88B491DE1DA92728D985CFE7C241D14FC15FDC5ACDA5B;
defparam prom_inst_3.INIT_RAM_11 = 256'h94049E51363CDA08C9A59EDCBBC4A651549267C822818F6E85CDD24A9104EDAE;
defparam prom_inst_3.INIT_RAM_12 = 256'h94D1561E6CA039241971075FE937CEB718C07D0DA1ED9D01523A600157959697;
defparam prom_inst_3.INIT_RAM_13 = 256'h0B5ADBBC0656AAB776901AEBB0447E13F05B59E3DF6568DF73E7F731C4AE23BF;
defparam prom_inst_3.INIT_RAM_14 = 256'h7E59ACE0F870E58CD2C41FFAC5631E64912944B2CEFAAED49EC3F716A88A4F02;
defparam prom_inst_3.INIT_RAM_15 = 256'h6CFC67803F001F8F77013AA7C963F0E076072D2F6B0932B270786F801DAABEBE;
defparam prom_inst_3.INIT_RAM_16 = 256'h007FFFFFFFFF800BFF4E9F87F0003235FFF03C1FFF8C61FFE0005FFE07038031;
defparam prom_inst_3.INIT_RAM_17 = 256'h2AA6084FEE57AF331FF6196C61775CBEEDFE3C363B388612790800100007FFFF;
defparam prom_inst_3.INIT_RAM_18 = 256'hD88B757731BE7145CADE2DCDD371CC6F2334C6175C4FF1A9C13DA8AD4E1276F8;
defparam prom_inst_3.INIT_RAM_19 = 256'h817F965C37022D5B13DF7752A069C5C5A2933683EF737B053B070DF39A4F99C4;
defparam prom_inst_3.INIT_RAM_1A = 256'hC90CD8514BB13C50179134B534068033791572479AFC7ECE1048D44633B7C0D8;
defparam prom_inst_3.INIT_RAM_1B = 256'hEF005670BBA1EC3C02D5801DB12AD7DCD33D44C6FC772E78DE115B41F27FA64F;
defparam prom_inst_3.INIT_RAM_1C = 256'h1C41FEC54A7F0FF0935B01E1AB6A18C148A5FE0DE989F8833C05EAE494BE3F64;
defparam prom_inst_3.INIT_RAM_1D = 256'h21FFD8BF0FC000FE0FF7E06FF01F8000178383A13FFFFB0F03BFD319A00FF40F;
defparam prom_inst_3.INIT_RAM_1E = 256'h0000014F8D90000000001E948007E36400000002000006DFFFFC02CE84000000;
defparam prom_inst_3.INIT_RAM_1F = 256'h000020218482000000000000013002000000000010FB5F6C0000000965FDC800;
defparam prom_inst_3.INIT_RAM_20 = 256'hAF82D4A97B92C33CAAAE0C475F6B488444FCFF5401C80200001FFD0000001000;
defparam prom_inst_3.INIT_RAM_21 = 256'h83C6CDE0873C4400AFFF36A2CF63FBC7DF950694930769720115670FD85A22D6;
defparam prom_inst_3.INIT_RAM_22 = 256'h22AD8255FF0AF6CE4530E737054E4570461CD954B202BAC4B9DEB310CFF1C04E;
defparam prom_inst_3.INIT_RAM_23 = 256'hC31DAD15CD116FB85A6F7CAFB525C5A58701652FB5AF0D2280610D93372199AE;
defparam prom_inst_3.INIT_RAM_24 = 256'h128F22F2108B1D73DB73A233A7636DC67B7B3DA4DF302DF00DA918A202609203;
defparam prom_inst_3.INIT_RAM_25 = 256'h181CE01BB273A66A56E59CEA526E8C2E65685E2D6495BF91B7827A2A01D397AD;
defparam prom_inst_3.INIT_RAM_26 = 256'hA6963ACD5B77599A3A992D3F89028F17522077BFF0FCEAFC8AA5D85AB3006719;
defparam prom_inst_3.INIT_RAM_27 = 256'h89F8A4CFE95DC062CCC1A3E6A074EF6DBE3B735F98EE3A809B82C07C0DCB746F;
defparam prom_inst_3.INIT_RAM_28 = 256'hB6D118CF6CD6B574037FC1C33345B5DE31476FFEF3619227D5293322E8D25BBC;
defparam prom_inst_3.INIT_RAM_29 = 256'h9CA407D960542F221077EAB83FB29F5ACA1C4DAB4AA11A882557DA14F30967D1;
defparam prom_inst_3.INIT_RAM_2A = 256'h6901435FDF13C102BA1921DE6728CE4F9E5BD3843FAE8F6276DED7B7F8384A74;
defparam prom_inst_3.INIT_RAM_2B = 256'hC17A1B2A82586EB2318979C5A286C7AA4563AB48CCD6D87D9F14DB462AC84FD8;
defparam prom_inst_3.INIT_RAM_2C = 256'h29B98F92AB8E7FF4D7A08805051969A6E8411CB75CF942F010137F62EEEFFD48;
defparam prom_inst_3.INIT_RAM_2D = 256'h21101D4740418E7C237B2A9F534FD43FE58888B526819A10EBD37E1964A066C7;
defparam prom_inst_3.INIT_RAM_2E = 256'hF00E33DF9FE3E3E7DC0238082F1798EECE4BD8F758AEE1F2D4114593BEDD635B;
defparam prom_inst_3.INIT_RAM_2F = 256'h00BF717E2F8005FFFFD2BD0F0801F071F838F8BABF81F83C805656188DF001F1;
defparam prom_inst_3.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000001E79E10;
defparam prom_inst_3.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_4 (
    .DO({prom_inst_4_dout_w[30:0],prom_inst_4_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_4.READ_MODE = 1'b0;
defparam prom_inst_4.BIT_WIDTH = 1;
defparam prom_inst_4.RESET_MODE = "SYNC";
defparam prom_inst_4.INIT_RAM_00 = 256'h00000000000000000000000000000000000000000000000000000000000002B2;
defparam prom_inst_4.INIT_RAM_01 = 256'h0000000000000000000000000006D90B0706D9102C1C1B6404B1706D9112C5C0;
defparam prom_inst_4.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_20 = 256'h48A90B93ACD437FB5F20145A108FBE5BB2D4C76C7D0B078B003CF4683017FFC0;
defparam prom_inst_4.INIT_RAM_21 = 256'h4086E46C8A9FA6DF89C7393489971964DE985B8BABDCD446C3F156B5595003DA;
defparam prom_inst_4.INIT_RAM_22 = 256'hDF1AE6A31928248A08938B9E39E1F23CE1BEF6AAE147404473EC3CFEB4A04548;
defparam prom_inst_4.INIT_RAM_23 = 256'hE0BB2B79CAE1C1025655506436CAAF4B29C8FF31E546BB1AB3C3EA2EBB15FF7B;
defparam prom_inst_4.INIT_RAM_24 = 256'h8C91F1C07E070F8065B7F1F00F1E31FED53031E3C078CF79553F3367F80CABC7;
defparam prom_inst_4.INIT_RAM_25 = 256'hCE70FC07F07C0000E3181E00FE1F00FE189807E03F0E07FF8C9801E0FE0F07FF;
defparam prom_inst_4.INIT_RAM_26 = 256'hF817FC01F500FF1C7F81FFF03F0001E38FFE07FC0780001E31E7E05FC0F00001;
defparam prom_inst_4.INIT_RAM_27 = 256'h52FB803EC8FFE2BF095FE857FC61EF8BFF500FFFABF861FC07FFA00FF40BE18F;
defparam prom_inst_4.INIT_RAM_28 = 256'hDDB57A1D075515FDCF16B7A5E9020814FF5F3C05F7FA955002FD57CE0A87FFD7;
defparam prom_inst_4.INIT_RAM_29 = 256'h4F1FC60E69BE1954A71151253DD6D2578C3C910809E109588DD6B207C89FC082;
defparam prom_inst_4.INIT_RAM_2A = 256'h766F6E69AF96735B022374D4CEEB6155B8E6FCF55F50025893FC7313B86A766C;
defparam prom_inst_4.INIT_RAM_2B = 256'h92E6AAA4C72623F2551E0ACC16CC076592393981B557B019F024AB1DE4BECE06;
defparam prom_inst_4.INIT_RAM_2C = 256'h7EC0E3636F478F5CFF83BE673D66C3CADB47F801FCF6A6197DE54C33112A0257;
defparam prom_inst_4.INIT_RAM_2D = 256'hA980E7C001E658F2657AADE78E824F9A4C20EA36A60E1FC29E6920A3E6CADC78;
defparam prom_inst_4.INIT_RAM_2E = 256'h5530AC7F8E1A1F319FF32AFCA9C38C3F8E663036D51D49C38C101C319C1A9502;
defparam prom_inst_4.INIT_RAM_2F = 256'hE0195B5C98FF0E007C39E386AB036C7FC7000F18E3E259112C7FC6040F18CFFB;
defparam prom_inst_4.INIT_RAM_30 = 256'hF0781FE326031C001F87FC3C7DF248F9B8783E03FC38E01949FD98FC1E007C38;
defparam prom_inst_4.INIT_RAM_31 = 256'hFFFFF407F0078E3F0F801FFFF83F800319FF1E007F8FF83C0F8333839C007F17;
defparam prom_inst_4.INIT_RAM_32 = 256'hFFFFFFFFE0007FFF81FB1FFFFFFFF000FFFFC3E003FFFFFFF80BFFFFC78007E4;
defparam prom_inst_4.INIT_RAM_33 = 256'h0000AFFFFFFFFD0000000000FFFFFFFFFC0017FCC017FFFFFFFFFE003FFF80FF;
defparam prom_inst_4.INIT_RAM_34 = 256'hFDF5FF34417C8353807FF0E3806527F19C3FF81401000001BBFFFFFFF8000000;
defparam prom_inst_4.INIT_RAM_35 = 256'hE652E39BA1F000F4B3F2AD9F2D6CFF6DC692CFB493E4FF0E3E07180D1AFA8BF8;
defparam prom_inst_4.INIT_RAM_36 = 256'hFF81E0FF8398E3E3FFEFF803C3C3CCDC0387FFFFF03CE00C923C703FFFFC0CE7;
defparam prom_inst_4.INIT_RAM_37 = 256'h1C3E000007C7DF8C4CFE30FC0000178FFF1DD9FC73E000800F83F839C71F07FF;
defparam prom_inst_4.INIT_RAM_38 = 256'h8CC1070FF9A007E0FFF399878E07FF4007E3FFE3333F1E1F80005FC3FFC6663E;
defparam prom_inst_4.INIT_RAM_39 = 256'h5BBDD3DEF42FFB7802FE03E1C73CFE0FF73E801E1FF0E6600F03FFFC0FF07FC3;
defparam prom_inst_4.INIT_RAM_3A = 256'hE7514F265D2EEC8E282E6F917715D46C31907530A2067A6B024AAF2D8E74BD54;
defparam prom_inst_4.INIT_RAM_3B = 256'h88C07E5AE794EDCCF9C84E6380ACD3DA0C0A59B92630D6CEB898BCA8D6130151;
defparam prom_inst_4.INIT_RAM_3C = 256'h0393003F0071F83807F1BB000FE0C1FFD87E0079B306B1FC07C03F078AD38E78;
defparam prom_inst_4.INIT_RAM_3D = 256'hFFE700400FF293CF381F1E00380F1C987F1E0E0FC0001F8327013E0F07F0A060;
defparam prom_inst_4.INIT_RAM_3E = 256'hF5099D2F7F599C67C090162A99D5A7C63CFEF8CA5157AB980300080386549E4C;
defparam prom_inst_4.INIT_RAM_3F = 256'h2F7B4566F620C4E14BB99B6682798C735FE66C6508EFA7E8686511031E960619;

pROM prom_inst_5 (
    .DO({prom_inst_5_dout_w[30:0],prom_inst_5_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_5.READ_MODE = 1'b0;
defparam prom_inst_5.BIT_WIDTH = 1;
defparam prom_inst_5.RESET_MODE = "SYNC";
defparam prom_inst_5.INIT_RAM_00 = 256'hC49A1D0B13DB673C85B0970A7AE365B9F2D77264FA411413E5398D46FAA09A31;
defparam prom_inst_5.INIT_RAM_01 = 256'h90FB1CD9D253605723A968E745E98ADD4D9D1AFBD225A43DB1419289687532C0;
defparam prom_inst_5.INIT_RAM_02 = 256'h564004C19B3191374EA1F0CE309669D4BA4467DCC4474E4182C3175084C779D2;
defparam prom_inst_5.INIT_RAM_03 = 256'h2A078BCB46CE253EFF746FAABA8028CD50D4E6222FAC9402954F70D41FBC8E56;
defparam prom_inst_5.INIT_RAM_04 = 256'hF625043A1DCADDB4A2CB562E120E7697E5AA344228ABCACC436B71E6A3D0D191;
defparam prom_inst_5.INIT_RAM_05 = 256'h1DC7272A64C3C94B0AC5F0B6A894FA57FA91867B1B44E96849E11804E7734110;
defparam prom_inst_5.INIT_RAM_06 = 256'hF7876DA13067C007E14C072DC5259FB3DB23F8210548F7AD27AC458ACF6B66B9;
defparam prom_inst_5.INIT_RAM_07 = 256'h8E4FE323FF800207FE1E1DEACE4C67F80100038FE1C65F272C00F8E040F1C981;
defparam prom_inst_5.INIT_RAM_08 = 256'hF03FC0077FFF2C007F0FF80FE03E03E000003F400783E70073C3F00007FFF247;
defparam prom_inst_5.INIT_RAM_09 = 256'h9ED41A9037FF00100000000001FFFFFFFFFC00003FF8007FFFFFFFFF800007FF;
defparam prom_inst_5.INIT_RAM_0A = 256'h09AF74FE960BD14824357C9F6C10ABEBA65960F645FF07F1C01101FDAE58A4C3;
defparam prom_inst_5.INIT_RAM_0B = 256'h67BEB369D30ED6DD1FE4EE314607BD25FEC9CDDB788FC8FA37243855DF9E297B;
defparam prom_inst_5.INIT_RAM_0C = 256'hFC3CA372024BE097731F5463F879458829B1F3CC042B0C07C99FAA00D8F5218C;
defparam prom_inst_5.INIT_RAM_0D = 256'h55547F1CC49DF11C1417AE82A4519E3C8EEC28B8CF1D668512F521E92E078382;
defparam prom_inst_5.INIT_RAM_0E = 256'h15C25F1C82921F374EA5A294C66D40039B7AC0AFD9B04B90B1390A949481DE2E;
defparam prom_inst_5.INIT_RAM_0F = 256'h727C1BB9F68F6276778A432BB08FA0383DC27177629FD1583E432957EA9F6A72;
defparam prom_inst_5.INIT_RAM_10 = 256'hB2FD8CAA7FC30DB63B07DA15B3FE077FCA009FBC45FF80E66BEA1475FF56A83A;
defparam prom_inst_5.INIT_RAM_11 = 256'hB3F8E00F6D1DD850A82CF0E0953FD6F6A3D5CC30C21CA5C29A4F11585601DB63;
defparam prom_inst_5.INIT_RAM_12 = 256'h068331FF8F0008006E591F4127080F48FBB60063AE80B31FA3C176D8B9E6E312;
defparam prom_inst_5.INIT_RAM_13 = 256'h7336387C0798F66D311A94F891C3FFE3800EC8E1D55B66230FFC78304D98D2EC;
defparam prom_inst_5.INIT_RAM_14 = 256'hAFCB63FF007F0045B10ACA36ACE01F871EE4AD83A25D85B3812319E99A59F2B7;
defparam prom_inst_5.INIT_RAM_15 = 256'h70FC1F803FFFFF80F0FE333838E000FF89FF1CE08DADCE6E0F806FFFFC667F2A;
defparam prom_inst_5.INIT_RAM_16 = 256'h007FFFFFFFFF800000B16007FFFFFFFFFFF003FFFFF07E001FFFFFFE00FF803E;
defparam prom_inst_5.INIT_RAM_17 = 256'h103610B1334BD2DAA7DC15CC6E0736CDA7EE4DD3BFF6E488D908001000000000;
defparam prom_inst_5.INIT_RAM_18 = 256'h93B84CD956E5DFF1D6FDD450B15F9F436D0AAF1AF330B7854C2D01C3058AC547;
defparam prom_inst_5.INIT_RAM_19 = 256'h0F76C15B1ECA382257D8A66474B64FC62690C5D61F18AD05623F823A2B117126;
defparam prom_inst_5.INIT_RAM_1A = 256'hE02067326CC3BE0C2F50EF65611AE10D0A8E98BC98967C80C80E250C9F07BF29;
defparam prom_inst_5.INIT_RAM_1B = 256'hE8A35A4672A67627BE655917DCDFA0EB0122F2DEAE06534703AD7B556F163DC1;
defparam prom_inst_5.INIT_RAM_1C = 256'h03C001067380FFF070C701FE324C07C73B9C000D8D2DFBB183FA1E6F7E78BFAB;
defparam prom_inst_5.INIT_RAM_1D = 256'h21FFFFFF003FFF000FFFFFFFF0007FFFE803FC5FFFFFFB00FFBFFC1E00000BFF;
defparam prom_inst_5.INIT_RAM_1E = 256'h0000014F8D90000000001E948007E36400000002000006DFFFFC000000000000;
defparam prom_inst_5.INIT_RAM_1F = 256'h000020218482000000000000013002000000000010FB5F6C0000000965FDC800;
defparam prom_inst_5.INIT_RAM_20 = 256'h8A41DFBA1842D210AB3AD5E3420018D1FFFC000400000200001FFD0000001000;
defparam prom_inst_5.INIT_RAM_21 = 256'hFBF316FF95F3683DDF62E48FB4A8FB51547406BA1FFEF603F1A376CC29B570F0;
defparam prom_inst_5.INIT_RAM_22 = 256'h82A88384D4FEBBF08D3C17372CD5EB3446C2AEE676AAAC9174EF64A305F957B4;
defparam prom_inst_5.INIT_RAM_23 = 256'h86D5E7053DB4C769EE7E6EAE3C627592F6624FE7648D3D372E96715486B43DF0;
defparam prom_inst_5.INIT_RAM_24 = 256'hB7B203F8A6F01CF0DBB0483F7B491B2574A6BB026F98956B02F76F6C1C804F5D;
defparam prom_inst_5.INIT_RAM_25 = 256'h88C3C412E3C4AE44EBA7A83331D074735FD624EF9D1DBAEFEDE3FF3AABD7432B;
defparam prom_inst_5.INIT_RAM_26 = 256'h2758C25B996064ECEF733704AD3CEB4D14F594099684C395C5DF6B99A289B0E0;
defparam prom_inst_5.INIT_RAM_27 = 256'hD2B5C95EB024E52A28A57A84E6DF94BF4A73DA2AE35B735203D86923687E04AF;
defparam prom_inst_5.INIT_RAM_28 = 256'hD1D7A6B38C28BC2381B5B2B8E07E3C77AF193B2936D39CB6314ABA1B228AD770;
defparam prom_inst_5.INIT_RAM_29 = 256'h88AF022A07599C99F95CC2B0EA8420E0B682DC317EF378B28BB8E20B6913DB50;
defparam prom_inst_5.INIT_RAM_2A = 256'hA418F7510B9BEA56E696149C139DE38D2B555B4A4E10A4F8B136F13256DB7CE0;
defparam prom_inst_5.INIT_RAM_2B = 256'h8AF3E8EA0CA2B72B61D9FE938EDD81004B3BC7DD7ADAC7FC46F9578D33B3E5D2;
defparam prom_inst_5.INIT_RAM_2C = 256'h1C55E2C1212DF2204855134857FA3885BAF71919888240640AB0A2DBB84FD0AC;
defparam prom_inst_5.INIT_RAM_2D = 256'h2330697296624191691CB301301683AD058A18736D86D3F4A886E0CEFB64EDAD;
defparam prom_inst_5.INIT_RAM_2E = 256'hF00FC3E0001FE0181FFE078FD94FD645C1C738F87FA10206521BD0707E331C6C;
defparam prom_inst_5.INIT_RAM_2F = 256'h00008E802FFFFFFFFFFFFD00F7FE007E07F800BFFF8007FC7F9B660783F0000F;
defparam prom_inst_5.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000001E79E10;
defparam prom_inst_5.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_5.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_6 (
    .DO({prom_inst_6_dout_w[30:0],prom_inst_6_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_6.READ_MODE = 1'b0;
defparam prom_inst_6.BIT_WIDTH = 1;
defparam prom_inst_6.RESET_MODE = "SYNC";
defparam prom_inst_6.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000002832;
defparam prom_inst_6.INIT_RAM_01 = 256'h0000000000000000000000000012B6489F12B600223C4AD84489F12B600223C0;
defparam prom_inst_6.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_20 = 256'hBB57D84863640C3388EA33C670F00183EE9879D3FEA5F9FF203FF07FBF57FFC0;
defparam prom_inst_6.INIT_RAM_21 = 256'h73520064467FCEDFD0AC9693A79607A06257F6869A183F34BEDC02733861FE13;
defparam prom_inst_6.INIT_RAM_22 = 256'h00FAF866154692740383FF7CACD74FC0981F11C2DB2CFF83E1F21E2E726FF938;
defparam prom_inst_6.INIT_RAM_23 = 256'hB70898FE0A933D57923330783347258E98C7FFC02CF7A2B6703FED8264B69AC8;
defparam prom_inst_6.INIT_RAM_24 = 256'hF0E1F03FFE00FF8079C7F00FFF01F000E63FF01FC007C08199C0F0E00003980A;
defparam prom_inst_6.INIT_RAM_25 = 256'h0F8003FFF003FFFF03E001FFFE00FFFFE0E0001FFF01FFFFF0E0001FFE00FFFF;
defparam prom_inst_6.INIT_RAM_26 = 256'h07FFFC000AFF001F807FFFF000FFFE03F001FFFC007FFFE03E001FFFC00FFFFE;
defparam prom_inst_6.INIT_RAM_27 = 256'h50057FC05F001FFF080017A8007E007FFF50000054007E03FFFFA0000BF401F0;
defparam prom_inst_6.INIT_RAM_28 = 256'h1E0007DD00000002301D405FE902000000A03FFABFFA95500002A80FF57FFFD7;
defparam prom_inst_6.INIT_RAM_29 = 256'hC70007FE187F9260DCD0002503C1016EAB268000081F01636B90E30280003FFD;
defparam prom_inst_6.INIT_RAM_2A = 256'h8780E6E63527F738FC3C0C4C33427D33870703CCC06523D670007CF0880CA478;
defparam prom_inst_6.INIT_RAM_2B = 256'h834B3A63C0D83C0E3303AD0C71C3F8780E77012C3D318FE1801D98E6B0CE467F;
defparam prom_inst_6.INIT_RAM_2C = 256'h7FFFE0EF0E90FECC0003BFFF0CE0EA8DC8C00001FFF19E1C51E33C00002FFE31;
defparam prom_inst_6.INIT_RAM_2D = 256'h987F07FFFFE1C7FCB6799C180FFFFF863C3AB3F261F01FFFFE18E0CA89D9C380;
defparam prom_inst_6.INIT_RAM_2E = 256'h99CF9C000FE5FF0F8003B303983C0FC07E1E0FC76603383C0FEFFC0F83E32601;
defparam prom_inst_6.INIT_RAM_2F = 256'hE01E63FC78000FFFFC07E00733FF1C0007FFFF07E00391EF1C0007FBFF07C003;
defparam prom_inst_6.INIT_RAM_30 = 256'hF007FFFC3800FC001FFFFC03FDFC70F878003FFFFC07E01E71FC78001FFFFC07;
defparam prom_inst_6.INIT_RAM_31 = 256'hFFFFF4000FF80FC0FF801FFFF8007FFC1E00FE007FFFF803FFFC3C007C007FFF;
defparam prom_inst_6.INIT_RAM_32 = 256'hFFFFFFFFE000000001FFFFFFFFFFF000000003FFFFFFFFFFF800000007FFFFE4;
defparam prom_inst_6.INIT_RAM_33 = 256'h0000AFFFFFFFFD0000000000FFFFFFFFFC0000000017FFFFFFFFFE00000000FF;
defparam prom_inst_6.INIT_RAM_34 = 256'hFFF5FF0DC1A900CF807FF01F8079C7F07C00001401000001BBFFFFFFF8000000;
defparam prom_inst_6.INIT_RAM_35 = 256'h079CFF87A1FFFFF38FFCC91F1CE3FF8E018E3FC6DC1C00FE01FF07F1ACF9B800;
defparam prom_inst_6.INIT_RAM_36 = 256'hFF801FFFFC1F001FFFFFF8003FC3F0E0007FFFFFF003E00F1C3C0FFFFFFC03E0;
defparam prom_inst_6.INIT_RAM_37 = 256'h03FE0000003FDFF070FE0FFC0000007FFFE1E1FC0FE00080007FFFC1F800FFFF;
defparam prom_inst_6.INIT_RAM_38 = 256'h0F0100FFF9A0001FFFFC1E0781FFFF40001FFFFC3C3F01FF8000003FFFF8783E;
defparam prom_inst_6.INIT_RAM_39 = 256'hC77DFC018BFFFB780001FFFE07C001FFF73E8001FFFF078000FFFFFC000FFFFC;
defparam prom_inst_6.INIT_RAM_3A = 256'hCAA8C0E2FD83CA6A6DE4D9F110E61D2458A1930F91F98198FC9320E07E0C022F;
defparam prom_inst_6.INIT_RAM_3B = 256'h783F81BA1FE6B1FBF8383FFC7C63669C43FA3B86381244BB2587F387DBDEAB97;
defparam prom_inst_6.INIT_RAM_3C = 256'hFC1C0000FFF007C7FFFE3C00001FC00027FFFF81C3FE0FFC003FFF000C9C01F8;
defparam prom_inst_6.INIT_RAM_3D = 256'hFFE0FFFFFFFCE3FF07FF01FFFFFFE0E07F01FE003FFFFFFC380101FF000F5F9F;
defparam prom_inst_6.INIT_RAM_3E = 256'h06077E353D387C1FC0EFF1CCD2339FC1FFFF07C06667987800FFFFFF8798E1C3;
defparam prom_inst_6.INIT_RAM_3F = 256'h9BA89AD4AD9F0DFE5CD7A03729F87DFC684E61B85A6F9FE7B0131E41D58E01F8;

pROM prom_inst_7 (
    .DO({prom_inst_7_dout_w[30:0],prom_inst_7_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_7.READ_MODE = 1'b0;
defparam prom_inst_7.BIT_WIDTH = 1;
defparam prom_inst_7.RESET_MODE = "SYNC";
defparam prom_inst_7.INIT_RAM_00 = 256'hBF8797C5A9426016FE8D693CA9A263EB8C4DEBD6A93E0C086354DAF4A99F09CF;
defparam prom_inst_7.INIT_RAM_01 = 256'hC684CA69C99C44501DA77F4AC30E73972D8C75134E8666E0B73D60825AC60CD2;
defparam prom_inst_7.INIT_RAM_02 = 256'hCF7AC9EAEABED502759E8A112BED669C448C1FCB6395B43BEE044D19D93A433E;
defparam prom_inst_7.INIT_RAM_03 = 256'hAB7D39526F7A3C7337F34FF3767FF0C33B99B99A9FB5B3FC8D85F40206140F71;
defparam prom_inst_7.INIT_RAM_04 = 256'h4F5EBE86BC34C66EEB82627266BED1B56D46324F8F84C59CEF3ACBBE7FE870E4;
defparam prom_inst_7.INIT_RAM_05 = 256'hFE4F1CE61FC3EF0F0DC75A7BD6CC2637E30DFE78250A4E73D8571806907F3A27;
defparam prom_inst_7.INIT_RAM_06 = 256'h0500E39FFF87C007E0CFF8C5C31C7FBC1F03FFE0C6BFEE631F9FC673CF0CE662;
defparam prom_inst_7.INIT_RAM_07 = 256'h0F8FE0E00000000001FFE1F33E3C18000100007FFE0760E0E3FF00E040F039FE;
defparam prom_inst_7.INIT_RAM_08 = 256'h003FFFFFFFFF2C0000F0000FFFC1FFE0000000BFF803F8000FC0000000000DB8;
defparam prom_inst_7.INIT_RAM_09 = 256'hEEAA23341BFF00100000000001FFFFFFFFFC00000000007FFFFFFFFF80000000;
defparam prom_inst_7.INIT_RAM_0A = 256'h536A78DCFF17FEAA93C67DB7F9471A68E1F800F87A00FFF1C01001FFBE51AFFF;
defparam prom_inst_7.INIT_RAM_0B = 256'h2430D90CA4A0A7456FB7BD4ADC37B3805495F4B0C1403B9D65D36891E39DBE56;
defparam prom_inst_7.INIT_RAM_0C = 256'h03FC800002481F687C1F43E0007FBF65EB8E211AE74CD8C822D6335F729FF80A;
defparam prom_inst_7.INIT_RAM_0D = 256'h8AF4006E727C3902C96FA00CC7BF83BC0013DF404F3A5BA412F5296181F803FD;
defparam prom_inst_7.INIT_RAM_0E = 256'h8C3C15B7C6721FB0C618CADB021D000078F2E437E38E40000F07F32723C6FE00;
defparam prom_inst_7.INIT_RAM_0F = 256'hCE0053FB067FFFF1CE344BF9047FFFFB8C3C5BBD067FFEFB8FBC43BD8E7F7FF1;
defparam prom_inst_7.INIT_RAM_10 = 256'hB56FCCB9FFFCFC71FB76DADA8FFFFF0E3A0ED6AEA3FFFFE31C8285F00CF6F7F9;
defparam prom_inst_7.INIT_RAM_11 = 256'h7000FFFF1CFDE37CEB9C00FF6F1C76EB6DF5DC00FDFC63C2EDB7D73817FFC71F;
defparam prom_inst_7.INIT_RAM_12 = 256'hE070F0000FFFF8E3FF9D910F1F000FFFF871FF8DE8878F0003FFF1C7FE3FE30E;
defparam prom_inst_7.INIT_RAM_13 = 256'h80F1F803F81F01E30FE327078FC00003FFFE381E199C9E1F00007FCFC387FCC8;
defparam prom_inst_7.INIT_RAM_14 = 256'h3038E000007FFFC38FF36C319C1FE007E01C6383349F9C707FFC1E0079C7FCDB;
defparam prom_inst_7.INIT_RAM_15 = 256'h7F03FF803FFFFF800FFFC3C007E000FFFFFF03E00E31FE1E00006FFFFC1E0033;
defparam prom_inst_7.INIT_RAM_16 = 256'h007FFFFFFFFF800000000007FFFFFFFFFFF0000000007FFFFFFFFFFE00007FC0;
defparam prom_inst_7.INIT_RAM_17 = 256'h2887CCDD68892D9179612274999B300D0C9F480B95E2A488D908001000000000;
defparam prom_inst_7.INIT_RAM_18 = 256'hB4D0A6D8C502CE9F966473F1EC493F3F004A466F48B609810184A6669ABB9FF2;
defparam prom_inst_7.INIT_RAM_19 = 256'h60CB8BEE0A6BDD4D3AC7947AC638ABE08C3D1535765FD4163C6FF56A4EACE651;
defparam prom_inst_7.INIT_RAM_1A = 256'h359FCECC9DA8B8C9AEB7EC20D3D3BA40E822A51001BC29F38AFECCF760BF7757;
defparam prom_inst_7.INIT_RAM_1B = 256'hEFDF36C0A9CA4D27C1D0B9B395D58108B350DDAD3507812ABC9D521CFC116871;
defparam prom_inst_7.INIT_RAM_1C = 256'h003FFFF87C00000FF03F01FFC38FFFC0F87C000DF1CE078F800001E3F8ACC767;
defparam prom_inst_7.INIT_RAM_1D = 256'h21FFFFFF000000000FFFFFFFF00000000003FFFFFFFFFB000040001FFFFFFFFF;
defparam prom_inst_7.INIT_RAM_1E = 256'h0000014F8D90000000001E948007E36400000002000006DFFFFC000000000000;
defparam prom_inst_7.INIT_RAM_1F = 256'h000020218482000000000000013002000000000010FB5F6C0000000965FDC800;
defparam prom_inst_7.INIT_RAM_20 = 256'h8001DFFA1002D210ABFE806352000AD4FFFC000400000200001FFD0000001000;
defparam prom_inst_7.INIT_RAM_21 = 256'h17C46DFF7566B37466DE1225868544CF2C0BF9401FFFFFFDF180880FF7F008FE;
defparam prom_inst_7.INIT_RAM_22 = 256'h7CB456C0306E6DBF0CEAB3B61C191D2C1348127C846D38376ECA93C6F9FB1D78;
defparam prom_inst_7.INIT_RAM_23 = 256'h1DF9BCFA037B8CE1DDBB1F4E1211A7318BC4B7E2CD5CDFEBC5F87CDD0FE81A3A;
defparam prom_inst_7.INIT_RAM_24 = 256'hA52DFB267F00F4B4CB2DDF68FC86BAF73C914E6FF00E8548F8CA751FE1E8BBCF;
defparam prom_inst_7.INIT_RAM_25 = 256'hB81DD749E387A59F5856A756F1E0C1CF8C2773BB7DE5B6651C0488EE6F8B6B8C;
defparam prom_inst_7.INIT_RAM_26 = 256'h35F5DD9DE72AD02C576E6CF8CEFA46002EFEE28618FC5A5427DE9548430F273E;
defparam prom_inst_7.INIT_RAM_27 = 256'h1CB3A4C0D537EC99EF39F9AD9F6D667AD9FC63F9A93BA92476B7F1BCE529069B;
defparam prom_inst_7.INIT_RAM_28 = 256'h702F8103F3E673C52DFC70781F87C3CD9F95CCD8F1CF9F380CD9BCA8444630FF;
defparam prom_inst_7.INIT_RAM_29 = 256'h837F0057F85FFC780198FFA7EA0000049EC1C3C26F1F07FA8000FDF8D8E29470;
defparam prom_inst_7.INIT_RAM_2A = 256'h63FFF0D01FFBD9310B5B3383FF83E3EE08CCD39068717FF80FF974CE31E5909F;
defparam prom_inst_7.INIT_RAM_2B = 256'hA60C081A60130289052F3A4F8EC3BF8FF0E95F9457063FFC3E019BFC967D66BE;
defparam prom_inst_7.INIT_RAM_2C = 256'hFF9E1E4FCC3C2740B0ECB6C06606E7C8CE25BE468A56C087F98F348292D27B95;
defparam prom_inst_7.INIT_RAM_2D = 256'hDF0F8E8E4E72880F18FFC3FF0FE7009B075F07F0E3871C0C68E4FDA40B3BE39C;
defparam prom_inst_7.INIT_RAM_2E = 256'h0FF003FFFFFFE0001FFE000FF8C01887C03F07007FA003FE31E261F001F0FF8F;
defparam prom_inst_7.INIT_RAM_2F = 256'h000000002FFFFFFFFFFFFD000000007FFFF800BFFF800003FFE386007FF00000;
defparam prom_inst_7.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000001E79E10;
defparam prom_inst_7.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_7.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_8 (
    .DO({prom_inst_8_dout_w[30:0],prom_inst_8_dout[4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_8.READ_MODE = 1'b0;
defparam prom_inst_8.BIT_WIDTH = 1;
defparam prom_inst_8.RESET_MODE = "SYNC";
defparam prom_inst_8.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000001575;
defparam prom_inst_8.INIT_RAM_01 = 256'h00000000000000000000000000DBB04CC7DBB039331F6EC0A0CD7DBB030335C8;
defparam prom_inst_8.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_20 = 256'hF91238381F8403C3FA3BF03E0F000003E11F803FFF9E01F8C03FF07FB097FFC0;
defparam prom_inst_8.INIT_RAM_21 = 256'h83CE0A9C3E000E201F9C34706068001F7E31218185E000F8FE448E0F078001E3;
defparam prom_inst_8.INIT_RAM_22 = 256'h0005001E18718E00007C00FF0E30C00087E00FF4871C00001E01FF49F1E00107;
defparam prom_inst_8.INIT_RAM_23 = 256'hC7F878000A8F019BEE0F0F8030C036F187C000001C04FC71F0001001E0DF0638;
defparam prom_inst_8.INIT_RAM_24 = 256'h00FE0FFFFE00007F81F80FFFFF000FFF07C00FFFC0003FFE1E000FE00000780C;
defparam prom_inst_8.INIT_RAM_25 = 256'h0FFFFFFFF000000003FFFFFFFE00000000FFFFFFFF00000000FFFFFFFE000000;
defparam prom_inst_8.INIT_RAM_26 = 256'hFFFFFC000000001FFFFFFFF000000003FFFFFFFC000000003FFFFFFFC0000000;
defparam prom_inst_8.INIT_RAM_27 = 256'h500000005FFFFFFF08000000007FFFFFFF50000000007FFFFFFFA000000001FF;
defparam prom_inst_8.INIT_RAM_28 = 256'h1FFFFFDD00000000001FFFFFE902000000003FFFFFFA95500000000FFFFFFFD7;
defparam prom_inst_8.INIT_RAM_29 = 256'h3F0007FE07FFE38083D00025003FFC7800DE80000800FE83D46FF30280000000;
defparam prom_inst_8.INIT_RAM_2A = 256'h07FFE1E039C7F0F8003FFC3C038C7D0F8007FFC3C079C3D1F0007FF0780F3878;
defparam prom_inst_8.INIT_RAM_2B = 256'h838C3A1FC0003FFE0F03CE0C0FC0007FFE0F01CE3D0F8001FFFC780738FE3E00;
defparam prom_inst_8.INIT_RAM_2C = 256'h7FFFE01F0F18FE3C0003BFFF03E0F30FC7C00001FFF07E1E61E0FC00002FFE0F;
defparam prom_inst_8.INIT_RAM_2D = 256'h780007FFFFE03FFF38787C000FFFFF81FC3CC3F1E0001FFFFE07E0F30FC7C000;
defparam prom_inst_8.INIT_RAM_2E = 256'h1E007C000FFFFF007FFC3C0078000FFFFE01FFF87800F8000FFFFC007FFC3800;
defparam prom_inst_8.INIT_RAM_2F = 256'h1FE07C03F8000FFFFC001FF83C00FC0007FFFF001FFC1E00FC0007FFFF003FFC;
defparam prom_inst_8.INIT_RAM_30 = 256'hF00000003FFFFC001FFFFC0002007F07F8003FFFFC001FE07E03F8001FFFFC00;
defparam prom_inst_8.INIT_RAM_31 = 256'hFFFFF40000000FFFFF801FFFF80000001FFFFE007FFFF80000003FFFFC007FFF;
defparam prom_inst_8.INIT_RAM_32 = 256'hFFFFFFFFE000000001FFFFFFFFFFF000000003FFFFFFFFFFF800000007FFFFE4;
defparam prom_inst_8.INIT_RAM_33 = 256'h0000AFFFFFFFFD0000000000FFFFFFFFFC0000000017FFFFFFFFFE00000000FF;
defparam prom_inst_8.INIT_RAM_34 = 256'hFFF5FF03C1CE003F807FF0007F81F80FFC00001401000001BBFFFFFFF8000000;
defparam prom_inst_8.INIT_RAM_35 = 256'hF81F007FA1FFFFF07FFF0E1F03E0000FFF81FFF8E003FFFE0000FFFE30F87800;
defparam prom_inst_8.INIT_RAM_36 = 256'hFF800000001FFFFFFFFFF800003C00FFFFFFFFFFF0001FF01FC3FFFFFFFC001F;
defparam prom_inst_8.INIT_RAM_37 = 256'hFFFE0000000020007F01FFFC000000000001FE03FFE0008000000001FFFFFFFF;
defparam prom_inst_8.INIT_RAM_38 = 256'h0FFEFFFFF9A0000000001FF87FFFFF40000000003FC0FFFF8000000000007FC1;
defparam prom_inst_8.INIT_RAM_39 = 256'hC0E2FFFFFFFFFB780000000007FFFFFFF73E8000000007FFFFFFFFFC00000000;
defparam prom_inst_8.INIT_RAM_3A = 256'h73983FE1FDC3262C463DC7F10FF81CE39D3E70FF80000007FF1C201FFE03C00F;
defparam prom_inst_8.INIT_RAM_3B = 256'hF8000005FFF8C1F807F8000003E07B1FC005F87FC00E38D3C3800F9FDC1E67E5;
defparam prom_inst_8.INIT_RAM_3C = 256'h001FFFFFFFF0000000003FFFFFFFC00000000001FC01FFFC000000FFF0E00007;
defparam prom_inst_8.INIT_RAM_3D = 256'hFFE000000000FC00FFFF0000000000FF80FFFE00000000003FFEFFFF00000000;
defparam prom_inst_8.INIT_RAM_3E = 256'hF800FFC64307FC003F000FF0E3F07FC00000003F878787F800000000781F003F;
defparam prom_inst_8.INIT_RAM_3F = 256'hD367BDDA638003FF904F9D1967F803FF8FDE616F39EF801FC00F1F95CC7E0007;

pROM prom_inst_9 (
    .DO({prom_inst_9_dout_w[30:0],prom_inst_9_dout[4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_9.READ_MODE = 1'b0;
defparam prom_inst_9.BIT_WIDTH = 1;
defparam prom_inst_9.RESET_MODE = "SYNC";
defparam prom_inst_9.INIT_RAM_00 = 256'h287ECBD3673C600D287CA312679C6018283CA1DA670003F84B33BDDA678007FF;
defparam prom_inst_9.INIT_RAM_01 = 256'hE33079D9C7E07D25FE7404D9C0F003B1B27910893E7818EB18FC58A6C63800C9;
defparam prom_inst_9.INIT_RAM_02 = 256'hC079F00C5B3F3880D380F9E0CC5E60F643A3FFC7801B7802480AC31FBE03A85E;
defparam prom_inst_9.INIT_RAM_03 = 256'h851C873C6079C3A17804FC090E0000C0FD0BC0271F6C70008203A544045A02CF;
defparam prom_inst_9.INIT_RAM_04 = 256'h80748D8183F8C7E0E4F981BF107E3076627E319170779B83DF1B783E000FCF07;
defparam prom_inst_9.INIT_RAM_05 = 256'h0035FC1E003C0F0F0FC73C03BA3C1E081C01FE783CF18EF63830E7F8F07F03EF;
defparam prom_inst_9.INIT_RAM_06 = 256'h06001F800007C007E0300009C0FC00401F03FFE038000BE0FF803803CF0FE61C;
defparam prom_inst_9.INIT_RAM_07 = 256'h0FF01FE000000000000001FC01FC0000010000000007801FE00000E040F00600;
defparam prom_inst_9.INIT_RAM_08 = 256'h003FFFFFFFFF2C000000000FFFFFFFE0000000000003FFFFFFC0000000000000;
defparam prom_inst_9.INIT_RAM_09 = 256'hFEE001B013FF00100000000001FFFFFFFFFC00000000007FFFFFFFFF80000000;
defparam prom_inst_9.INIT_RAM_0A = 256'h3713A0CA405579998FF87C700E67FA17E007FF007FFFFFF1C01001FFBE51AFFF;
defparam prom_inst_9.INIT_RAM_0B = 256'h56FDB70EC79A686E3C92606CBD6C4528B24C06DFD4BF5113134FB2ECA86910B1;
defparam prom_inst_9.INIT_RAM_0C = 256'hFFFC8000024800007FE0BFE0007FFF1C15C8CCC618703A203465293F9CFC9473;
defparam prom_inst_9.INIT_RAM_0D = 256'h000BFF8F8003F90000005FF0F8007FBC000000004F3FFFA412F52060000003FF;
defparam prom_inst_9.INIT_RAM_0E = 256'h7C00663B41F21FB03E00F31FC1FD000007F2F8C7E07E400000FFFC38003FFE00;
defparam prom_inst_9.INIT_RAM_0F = 256'h3E00623FC1FFFFF03E00723FC3FFFFF87C00623BC1FFFFF87E00723B49FF7FF0;
defparam prom_inst_9.INIT_RAM_10 = 256'hB78E0C87FFFFFC0FFB78E2D87FFFFF01FA0F18BE1FFFFFE0FC82E67D83F6FFF8;
defparam prom_inst_9.INIT_RAM_11 = 256'hF000FFFF03FDFC60E87C00FFFF03F6FC71F43C00FFFC1FC2F1C7D0F817FFC0FF;
defparam prom_inst_9.INIT_RAM_12 = 256'h000FF0000FFFF81FFFE1E100FF000FFFF80FFFF1D0807F0003FFF03FFFC70301;
defparam prom_inst_9.INIT_RAM_13 = 256'h000FF800001FFFE0FFFC38007FC00003FFFE07FFE1E001FF00007FFFC07FFF0F;
defparam prom_inst_9.INIT_RAM_14 = 256'hC007E000007FFFC07FFC70307C000007FFFC1F83C71F83F000001FFFF83FFF1C;
defparam prom_inst_9.INIT_RAM_15 = 256'h7FFFFF803FFFFF80000003FFFFE000FFFFFF001FF03E01FE00006FFFFC01FFC3;
defparam prom_inst_9.INIT_RAM_16 = 256'h007FFFFFFFFF800000000007FFFFFFFFFFF0000000007FFFFFFFFFFE00000000;
defparam prom_inst_9.INIT_RAM_17 = 256'h3DDE7A600A482AF96B7F920E234899D4E187291E03B2A488D908001000000000;
defparam prom_inst_9.INIT_RAM_18 = 256'hD808A67EA740C06897FAD902C454598A6DB5E52C593FC9593DAD7B96E3C12DD4;
defparam prom_inst_9.INIT_RAM_19 = 256'hCC8EDCCC0A4ADD4C4AD7B672A4288D966633B966630ECE606F5366737EB37E77;
defparam prom_inst_9.INIT_RAM_1A = 256'hB7CC21FFFC67BF6DC87013E3CFDCCC7FE801630FE339A00CFB320000009FFFDD;
defparam prom_inst_9.INIT_RAM_1B = 256'hEFFF0E3F32F1A327FFCC79DAE43381F788C0960A1307FF1980D79E33FFEF1BC1;
defparam prom_inst_9.INIT_RAM_1C = 256'h000000007FFFFFFFF000FE0003F0003FF803FFF201F0007F8000001FFF30FF1F;
defparam prom_inst_9.INIT_RAM_1D = 256'h21FFFFFF000000000FFFFFFFF00000000003FFFFFFFFFB000000001FFFFFFFFF;
defparam prom_inst_9.INIT_RAM_1E = 256'h0000014F8D90000000001E948007E36400000002000006DFFFFC000000000000;
defparam prom_inst_9.INIT_RAM_1F = 256'h000020218482000000000000013002000000000010FB5F6C0000000965FDC800;
defparam prom_inst_9.INIT_RAM_20 = 256'h8001DFFA1002D210ABFE8263520008D4FFFC000400000200001FFD0000001000;
defparam prom_inst_9.INIT_RAM_21 = 256'hA61C23FFF4EE0255663E0E6387367FC0FC0000001FFFFFFFF180000FFFF000FE;
defparam prom_inst_9.INIT_RAM_22 = 256'hFF43CE437C03847FF3E6703C61A4FEC3CEC714C78DEFC78CE0E38511FE073300;
defparam prom_inst_9.INIT_RAM_23 = 256'h5A1A63FFFF084C95A186FFF1F1098ABC34BCF81E2301CF0E23FF83CC80F8C349;
defparam prom_inst_9.INIT_RAM_24 = 256'h2AEF0E11FFFFF38CCC7A18E7FFFF861721E8611FFFFE72C88B430CFFFFE787C8;
defparam prom_inst_9.INIT_RAM_25 = 256'h8F5A10C7E3F85C4243A54C31F1FF3C2101D68618FDFA4E2301D60E19EFFCF852;
defparam prom_inst_9.INIT_RAM_26 = 256'hC433C01E00E6303168611C00F0062101D78611801F03C6343AF0C33803F0D084;
defparam prom_inst_9.INIT_RAM_27 = 256'h1F4F9C3F19B81C78103E079C7F89B80638007C0798FBCDB80E7001C01CE7072D;
defparam prom_inst_9.INIT_RAM_28 = 256'h0FFF8003FFE1F00631FC0FF80007FFC380198FF80FC0603FFC3840CC7FC1F000;
defparam prom_inst_9.INIT_RAM_29 = 256'h7FFF0000005FFC07FE1F005FEA0000009EC03FFC7000FFFA8000FFF838031870;
defparam prom_inst_9.INIT_RAM_2A = 256'h1FFFF02FE3E438F00C63307FFF801C0FF7C3D3E3880FFFF8000077FE0FFE1F00;
defparam prom_inst_9.INIT_RAM_2B = 256'h9E000805FF1C0198F9B2C63F8EC07FF38018C0199FC1FFFC01FE1C038E0188FE;
defparam prom_inst_9.INIT_RAM_2C = 256'h001FFE3FF1CC113F45C38E3F87FE1FF10E137FA569CE3F07F87FC702763C5D63;
defparam prom_inst_9.INIT_RAM_2D = 256'hFF000FFE3E7CF000F80003FF0007FF870610000FE0781FFC1707039C0C43E07C;
defparam prom_inst_9.INIT_RAM_2E = 256'h000003FFFFFFE0001FFE000FF83FE0F83FFF00007FA003FE0FFC7E0FFFF0000F;
defparam prom_inst_9.INIT_RAM_2F = 256'h000000002FFFFFFFFFFFFD000000007FFFF800BFFF8000000003F9FFFFF00000;
defparam prom_inst_9.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000001E79E10;
defparam prom_inst_9.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_9.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_10 (
    .DO({prom_inst_10_dout_w[30:0],prom_inst_10_dout[5]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_10.READ_MODE = 1'b0;
defparam prom_inst_10.BIT_WIDTH = 1;
defparam prom_inst_10.RESET_MODE = "SYNC";
defparam prom_inst_10.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000000033;
defparam prom_inst_10.INIT_RAM_01 = 256'h0000000000000000000000000092B0580792B08C605E4AC21581792B09C601E5;
defparam prom_inst_10.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_20 = 256'hF8E407F800040003F9CC0FFE00000003E01FFFFFFF8001F8003FF07FB017FFC0;
defparam prom_inst_10.INIT_RAM_21 = 256'h03C1F303FE000E001F83D80FE00000007E0E407F80000000FE3901FF00000003;
defparam prom_inst_10.INIT_RAM_22 = 256'h00000001E1807E0000000000300FC0008000000700FC0000000000700FE00100;
defparam prom_inst_10.INIT_RAM_23 = 256'hF807F8000A80FE1C01FF0000303FC7007FC0000003F8C00FF00000001F1801F8;
defparam prom_inst_10.INIT_RAM_24 = 256'h00FFFFFFFE00000001FFFFFFFF00000007FFFFFFC00000001FFFFFE0000007F0;
defparam prom_inst_10.INIT_RAM_25 = 256'h0FFFFFFFF000000003FFFFFFFE00000000FFFFFFFF00000000FFFFFFFE000000;
defparam prom_inst_10.INIT_RAM_26 = 256'hFFFFFC000000001FFFFFFFF000000003FFFFFFFC000000003FFFFFFFC0000000;
defparam prom_inst_10.INIT_RAM_27 = 256'h500000005FFFFFFF08000000007FFFFFFF50000000007FFFFFFFA000000001FF;
defparam prom_inst_10.INIT_RAM_28 = 256'h1FFFFFDD00000000001FFFFFE902000000003FFFFFFA95500000000FFFFFFFD7;
defparam prom_inst_10.INIT_RAM_29 = 256'hFF0007FE000003FF7FD000250000007FFFFE800008000003FFFFF30280000000;
defparam prom_inst_10.INIT_RAM_2A = 256'h07FFE01FC1F80FF8003FFC03FC0F82FF8007FFC03F81FC2FF0007FF007F03F87;
defparam prom_inst_10.INIT_RAM_2B = 256'h7C0FC5FFC0003FFE00FC0FF3FFC0007FFE00FE0FC2FF8001FFFC07F83F01FE00;
defparam prom_inst_10.INIT_RAM_2C = 256'h7FFFE000F01F01FC0003BFFF001F03F03FC00001FFF001E07E1FFC00002FFE00;
defparam prom_inst_10.INIT_RAM_2D = 256'hF80007FFFFE000003F87FC000FFFFF8003C0FC0FE0001FFFFE001F03F03FC000;
defparam prom_inst_10.INIT_RAM_2E = 256'h1FFFFC000FFFFF0000003FFFF8000FFFFE0000007FFFF8000FFFFC0000003FFF;
defparam prom_inst_10.INIT_RAM_2F = 256'h00007FFFF8000FFFFC0000003FFFFC0007FFFF0000001FFFFC0007FFFF000000;
defparam prom_inst_10.INIT_RAM_30 = 256'hF00000003FFFFC001FFFFC0000007FFFF8003FFFFC0000007FFFF8001FFFFC00;
defparam prom_inst_10.INIT_RAM_31 = 256'hFFFFF40000000FFFFF801FFFF80000001FFFFE007FFFF80000003FFFFC007FFF;
defparam prom_inst_10.INIT_RAM_32 = 256'hFFFFFFFFE000000001FFFFFFFFFFF000000003FFFFFFFFFFF800000007FFFFE4;
defparam prom_inst_10.INIT_RAM_33 = 256'h0000AFFFFFFFFD0000000000FFFFFFFFFC0000000017FFFFFFFFFE00000000FF;
defparam prom_inst_10.INIT_RAM_34 = 256'hFFF5FF003E0FFFFF807FF0000001FFFFFC00001401000001BBFFFFFFF8000000;
defparam prom_inst_10.INIT_RAM_35 = 256'h001FFFFFA1FFFFF000000FE0FFE0000FFF800000FFFFFFFE000000003F07F800;
defparam prom_inst_10.INIT_RAM_36 = 256'hFF800000001FFFFFFFFFF800000000FFFFFFFFFFF00000001FFFFFFFFFFC0000;
defparam prom_inst_10.INIT_RAM_37 = 256'hFFFE0000000000007FFFFFFC000000000001FFFFFFE0008000000001FFFFFFFF;
defparam prom_inst_10.INIT_RAM_38 = 256'h0FFFFFFFF9A0000000001FFFFFFFFF40000000003FFFFFFF8000000000007FFF;
defparam prom_inst_10.INIT_RAM_39 = 256'hC000FFFFFFFFFB780000000007FFFFFFF73E8000000007FFFFFFFFFC00000000;
defparam prom_inst_10.INIT_RAM_3A = 256'h8387FFE00203E1EF883C3FF100001C1FE1C00FFF80000000001FDFFFFE00000F;
defparam prom_inst_10.INIT_RAM_3B = 256'hF80000000000FE07FFF80000001F83E03FFFF8000001FF1C007FFF80201E1FF9;
defparam prom_inst_10.INIT_RAM_3C = 256'h001FFFFFFFF0000000003FFFFFFFC00000000001FFFFFFFC0000000000FFFFFF;
defparam prom_inst_10.INIT_RAM_3D = 256'hFFE000000000FFFFFFFF0000000000FFFFFFFE00000000003FFFFFFF00000000;
defparam prom_inst_10.INIT_RAM_3E = 256'h0000000780FFFC0000000000FC0FFFC00000000007F87FF800000000001FFFFF;
defparam prom_inst_10.INIT_RAM_3F = 256'h1CE07E9E1F8000001FC07E5F1FF800000FC19E4F07EF80000000E019C3FE0000;

pROM prom_inst_11 (
    .DO({prom_inst_11_dout_w[30:0],prom_inst_11_dout[5]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_11.READ_MODE = 1'b0;
defparam prom_inst_11.BIT_WIDTH = 1;
defparam prom_inst_11.RESET_MODE = "SYNC";
defparam prom_inst_11.INIT_RAM_00 = 256'hCFFE429F1F006003CFFC625E1F806007CFFC629E1F0000078CF07E9E1F800000;
defparam prom_inst_11.INIT_RAM_01 = 256'hFE857839C0007CF9FFEC57C7C000038E3FFB1AF8FE0000E7DFFCC23E3E0000C7;
defparam prom_inst_11.INIT_RAM_02 = 256'hC078000FC43FF42BCF80F8000FC060F26B9FFFC0001F0003D8AE3F1F8003E79E;
defparam prom_inst_11.INIT_RAM_03 = 256'h9E5C7F006078003F0007DEB8FE0000C001F8003E95E3F00080003B3807C8AE3F;
defparam prom_inst_11.INIT_RAM_04 = 256'h00732C7F8000C7E0E0F8003EE401F008607E301F0007BD003F04783E000FC007;
defparam prom_inst_11.INIT_RAM_05 = 256'h000603FE00000F0F0FC700038303FE000001FE783C000E0407F00000F07F03E0;
defparam prom_inst_11.INIT_RAM_06 = 256'h07FFFF800007C007E000000E3FFC00001F03FFE000000C1FFF800003CF0FE600;
defparam prom_inst_11.INIT_RAM_07 = 256'h0FFFFFE000000000000001FFFFFC0000010000000007FFFFE00000E040F00000;
defparam prom_inst_11.INIT_RAM_08 = 256'h003FFFFFFFFF2C000000000FFFFFFFE0000000000003FFFFFFC0000000000000;
defparam prom_inst_11.INIT_RAM_09 = 256'hFEE0003003FF00100000000001FFFFFFFFFC00000000007FFFFFFFFF80000000;
defparam prom_inst_11.INIT_RAM_0A = 256'hF0FC3F39C0667F8780007C0FF07805FFE00000007FFFFFF1C01001FFBE51AFFF;
defparam prom_inst_11.INIT_RAM_0B = 256'h98FC70F0F879E077BF8E1F8F031C0630F1C3F8E03380621F0F3FC303980E20F0;
defparam prom_inst_11.INIT_RAM_0C = 256'hFFFC8000024800007FFFFFE0007FFF03FE0F003E007FF9E0388727001F038C03;
defparam prom_inst_11.INIT_RAM_0D = 256'h0000000FFFFFF90000000000FFFFFFBC000000004F3FFFA412F52060000003FF;
defparam prom_inst_11.INIT_RAM_0E = 256'h03FF87C03FF21FB001FF03E03FFD0000000D00F81FFE40000000003FFFFFFE00;
defparam prom_inst_11.INIT_RAM_0F = 256'h01FF83C03FFFFFF001FF83C03FFFFFF803FF83C03FFFFFF801FF83C037FF7FF0;
defparam prom_inst_11.INIT_RAM_10 = 256'h480FF37FFFFFFC000480FD27FFFFFF0005F01F41FFFFFFE0037D07827FF6FFF8;
defparam prom_inst_11.INIT_RAM_11 = 256'hF000FFFF0002007F17FC00FFFF0009007E0BFC00FFFC003D01F82FF817FFC000;
defparam prom_inst_11.INIT_RAM_12 = 256'hFFFFF0000FFFF8000001FEFFFF000FFFF8000001FF7FFF0003FFF0000007FCFF;
defparam prom_inst_11.INIT_RAM_13 = 256'hFFFFF800001FFFE000003FFFFFC00003FFFE000001FFFFFF00007FFFC000000F;
defparam prom_inst_11.INIT_RAM_14 = 256'hFFFFE000007FFFC000007FCFFC000007FFFC007C07E07FF000001FFFF800001F;
defparam prom_inst_11.INIT_RAM_15 = 256'h7FFFFF803FFFFF80000003FFFFE000FFFFFF0000003FFFFE00006FFFFC000003;
defparam prom_inst_11.INIT_RAM_16 = 256'h007FFFFFFFFF800000000007FFFFFFFFFFF0000000007FFFFFFFFFFE00000000;
defparam prom_inst_11.INIT_RAM_17 = 256'hACCE6A644A492AD96B76924FA54A54CCC997291B13B2A488D908001000000000;
defparam prom_inst_11.INIT_RAM_18 = 256'hD448A6766A74C95996ECD991A454F1819999A52D5936A5492AA00C0C137A7881;
defparam prom_inst_11.INIT_RAM_19 = 256'hCCCECCCC0A4ADD4C4AD7B672A4288DCCCC999966664ECC446E6766733B337666;
defparam prom_inst_11.INIT_RAM_1A = 256'hC60C1FFFFC1FBF8E080FFFE03FDF0F8017FFE0FFFC3FDFFFFB320000009FFFDD;
defparam prom_inst_11.INIT_RAM_1B = 256'hEFFF01FFC3001F27FFC3F9E3040F81FF87C0E70E0F07FF0780E61E0FFFFF07C1;
defparam prom_inst_11.INIT_RAM_1C = 256'h000000007FFFFFFFF000000003FFFFFFF800000001FFFFFF80000000003F00FF;
defparam prom_inst_11.INIT_RAM_1D = 256'h21FFFFFF000000000FFFFFFFF00000000003FFFFFFFFFB000000001FFFFFFFFF;
defparam prom_inst_11.INIT_RAM_1E = 256'h0000014F8D90000000001E948007E36400000002000006DFFFFC000000000000;
defparam prom_inst_11.INIT_RAM_1F = 256'h000020218482000000000000013002000000000010FB5F6C0000000965FDC800;
defparam prom_inst_11.INIT_RAM_20 = 256'h8001DFFA1002D210ABFE8063520008D4FFFC000400000200001FFD0000001000;
defparam prom_inst_11.INIT_RAM_21 = 256'hC41C1FFFF41E039A6601FE1F87C7803FFC0000001FFFFFFFF180000FFFF000FE;
defparam prom_inst_11.INIT_RAM_22 = 256'hFFFFC1C0784383FFFFE1F0384183FFFFC1C0188783EFFF83E0F3070FFFFF0F00;
defparam prom_inst_11.INIT_RAM_23 = 256'h9C181FFFFF07CCF9C181FFFFF0F98F38307CFFFE1F01EE0E1FFFFFC380F08307;
defparam prom_inst_11.INIT_RAM_24 = 256'h23CE0E0FFFFFF07CCFBC181FFFFF81F73EF060FFFFFE0FC8F38303FFFFE07FCF;
defparam prom_inst_11.INIT_RAM_25 = 256'h8F9C103FE3FFFC3E43C60C0FF1FFFC1F01E70607FDFFFE1F01E70E07EFFFF83E;
defparam prom_inst_11.INIT_RAM_26 = 256'h040FC01FFFE1F03E7060FC00FFFE1F01E7060F801FFFC1F43CE0C0F803FFF07C;
defparam prom_inst_11.INIT_RAM_27 = 256'h1FFF83FFE1C003F8003FFF83FFF1C001F8007FFF87FBF1C001F001FFFC1F07CE;
defparam prom_inst_11.INIT_RAM_28 = 256'hFFFF8003FFE00FF83E03FFF80007FFC07FE1F007FFC0003FFC07FF0F803FF000;
defparam prom_inst_11.INIT_RAM_29 = 256'hFFFF0000005FFC00001FFFFFEA0000009EC000007FFFFFFA8000FFF807FC1F8F;
defparam prom_inst_11.INIT_RAM_2A = 256'hFFFFF00003FFF80FF07CCFFFFF80000FFFC02C03F7FFFFF8000077FE00001FFF;
defparam prom_inst_11.INIT_RAM_2B = 256'h7E000800001FFF87FE3C01FF8EC00003FFF83FE1E03FFFFC00001FFF81FE0F01;
defparam prom_inst_11.INIT_RAM_2C = 256'h001FFE0001F3F0FF86007E0007FE0001F1F0FFC6083E0007F80007FDF1FF9E00;
defparam prom_inst_11.INIT_RAM_2D = 256'hFF000FFE0180FFFFF80003FF0007FF80F81FFFFFE0001FFC0007FF83F07C1FFC;
defparam prom_inst_11.INIT_RAM_2E = 256'h000003FFFFFFE0001FFE000FF80000FFFFFF00007FA003FE00007FFFFFF0000F;
defparam prom_inst_11.INIT_RAM_2F = 256'h000000002FFFFFFFFFFFFD000000007FFFF800BFFF8000000003FFFFFFF00000;
defparam prom_inst_11.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000001E79E10;
defparam prom_inst_11.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_12 (
    .DO({prom_inst_12_dout_w[30:0],prom_inst_12_dout[6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_12.READ_MODE = 1'b0;
defparam prom_inst_12.BIT_WIDTH = 1;
defparam prom_inst_12.RESET_MODE = "SYNC";
defparam prom_inst_12.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000005545;
defparam prom_inst_12.INIT_RAM_01 = 256'h00000000000000000000000001B6B46A0FB6B491A87EDAD262A0FB6B488A83E0;
defparam prom_inst_12.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_12.INIT_RAM_20 = 256'hF807FFF800040003F80FFFFE00000003E01FFFFFFF8001F8003FF07FB017FFC0;
defparam prom_inst_12.INIT_RAM_21 = 256'h03C003FFFE000E001F801FFFE00000007E007FFF80000000FE01FFFF00000003;
defparam prom_inst_12.INIT_RAM_22 = 256'h0000000001FFFE00000000003FFFC00080000007FFFC00000000007FFFE00100;
defparam prom_inst_12.INIT_RAM_23 = 256'hFFFFF8000A80001FFFFF0000300007FFFFC000000000FFFFF0000000001FFFF8;
defparam prom_inst_12.INIT_RAM_24 = 256'h00FFFFFFFE00000001FFFFFFFF00000007FFFFFFC00000001FFFFFE000000000;
defparam prom_inst_12.INIT_RAM_25 = 256'h0FFFFFFFF000000003FFFFFFFE00000000FFFFFFFF00000000FFFFFFFE000000;
defparam prom_inst_12.INIT_RAM_26 = 256'hFFFFFC000000001FFFFFFFF000000003FFFFFFFC000000003FFFFFFFC0000000;
defparam prom_inst_12.INIT_RAM_27 = 256'h500000005FFFFFFF08000000007FFFFFFF50000000007FFFFFFFA000000001FF;
defparam prom_inst_12.INIT_RAM_28 = 256'h1FFFFFDD00000000001FFFFFE902000000003FFFFFFA95500000000FFFFFFFD7;
defparam prom_inst_12.INIT_RAM_29 = 256'hFF0007FE000003FFFFD000250000007FFFFE800008000003FFFFF30280000000;
defparam prom_inst_12.INIT_RAM_2A = 256'h07FFE00001FFFFF8003FFC00000FFFFF8007FFC00001FFFFF0007FF000003FFF;
defparam prom_inst_12.INIT_RAM_2B = 256'h000FFFFFC0003FFE00000FFFFFC0007FFE00000FFFFF8001FFFC00003FFFFE00;
defparam prom_inst_12.INIT_RAM_2C = 256'h7FFFE000001FFFFC0003BFFF000003FFFFC00001FFF000007FFFFC00002FFE00;
defparam prom_inst_12.INIT_RAM_2D = 256'hF80007FFFFE000003FFFFC000FFFFF800000FFFFE0001FFFFE000003FFFFC000;
defparam prom_inst_12.INIT_RAM_2E = 256'h1FFFFC000FFFFF0000003FFFF8000FFFFE0000007FFFF8000FFFFC0000003FFF;
defparam prom_inst_12.INIT_RAM_2F = 256'h00007FFFF8000FFFFC0000003FFFFC0007FFFF0000001FFFFC0007FFFF000000;
defparam prom_inst_12.INIT_RAM_30 = 256'hF00000003FFFFC001FFFFC0000007FFFF8003FFFFC0000007FFFF8001FFFFC00;
defparam prom_inst_12.INIT_RAM_31 = 256'hFFFFF40000000FFFFF801FFFF80000001FFFFE007FFFF80000003FFFFC007FFF;
defparam prom_inst_12.INIT_RAM_32 = 256'hFFFFFFFFE000000001FFFFFFFFFFF000000003FFFFFFFFFFF800000007FFFFE4;
defparam prom_inst_12.INIT_RAM_33 = 256'h0000AFFFFFFFFD0000000000FFFFFFFFFC0000000017FFFFFFFFFE00000000FF;
defparam prom_inst_12.INIT_RAM_34 = 256'hFFF5FF00000FFFFF807FF0000001FFFFFC00001401000001BBFFFFFFF8000000;
defparam prom_inst_12.INIT_RAM_35 = 256'h001FFFFFA1FFFFF000000FFFFFE0000FFF800000FFFFFFFE000000003FFFF800;
defparam prom_inst_12.INIT_RAM_36 = 256'hFF800000001FFFFFFFFFF800000000FFFFFFFFFFF00000001FFFFFFFFFFC0000;
defparam prom_inst_12.INIT_RAM_37 = 256'hFFFE0000000000007FFFFFFC000000000001FFFFFFE0008000000001FFFFFFFF;
defparam prom_inst_12.INIT_RAM_38 = 256'h0FFFFFFFF9A0000000001FFFFFFFFF40000000003FFFFFFF8000000000007FFF;
defparam prom_inst_12.INIT_RAM_39 = 256'hC000FFFFFFFFFB780000000007FFFFFFF73E8000000007FFFFFFFFFC00000000;
defparam prom_inst_12.INIT_RAM_3A = 256'hFC7FFFE00003E0100FC3FFF100001C0001FFFFFF80000000001FFFFFFE00000F;
defparam prom_inst_12.INIT_RAM_3B = 256'hF80000000000FFFFFFF80000000003FFFFFFF8000000001FFFFFFF80001E0001;
defparam prom_inst_12.INIT_RAM_3C = 256'h001FFFFFFFF0000000003FFFFFFFC00000000001FFFFFFFC0000000000FFFFFF;
defparam prom_inst_12.INIT_RAM_3D = 256'hFFE000000000FFFFFFFF0000000000FFFFFFFE00000000003FFFFFFF00000000;
defparam prom_inst_12.INIT_RAM_3E = 256'h00000007FFFFFC0000000000FFFFFFC00000000007FFFFF800000000001FFFFF;
defparam prom_inst_12.INIT_RAM_3F = 256'h1FE000E1FF8000001FC00060FFF800000FC00070FFEF80000000001E3FFE0000;

pROM prom_inst_13 (
    .DO({prom_inst_13_dout_w[30:0],prom_inst_13_dout[6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_13.READ_MODE = 1'b0;
defparam prom_inst_13.BIT_WIDTH = 1;
defparam prom_inst_13.RESET_MODE = "SYNC";
defparam prom_inst_13.INIT_RAM_00 = 256'h0FFE3CE0FF0060000FFC1C61FF8060000FFC1CE1FF0000000FF000E1FF800000;
defparam prom_inst_13.INIT_RAM_01 = 256'hFE7987F9C0007C01FFE3983FC00003803FF8E307FE0000E01FFC3CC1FE0000C0;
defparam prom_inst_13.INIT_RAM_02 = 256'hC078000FC03FF3CC3F80F8000FC060F18C7FFFC0001F0003C731FF1F8003E01E;
defparam prom_inst_13.INIT_RAM_03 = 256'h8063FF006078003F0007C0C7FE0000C001F8003E661FF00080003F0007C731FF;
defparam prom_inst_13.INIT_RAM_04 = 256'h007033FF8000C7E0E0F8003E07FFF000607E301F000781FFFF00783E000FC007;
defparam prom_inst_13.INIT_RAM_05 = 256'h0007FFFE00000F0F0FC7000383FFFE000001FE783C000E07FFF00000F07F03E0;
defparam prom_inst_13.INIT_RAM_06 = 256'h07FFFF800007C007E000000FFFFC00001F03FFE000000FFFFF800003CF0FE600;
defparam prom_inst_13.INIT_RAM_07 = 256'h0FFFFFE000000000000001FFFFFC0000010000000007FFFFE00000E040F00000;
defparam prom_inst_13.INIT_RAM_08 = 256'h003FFFFFFFFF2C000000000FFFFFFFE0000000000003FFFFFFC0000000000000;
defparam prom_inst_13.INIT_RAM_09 = 256'hFEE0003003FF00100000000001FFFFFFFFFC00000000007FFFFFFFFF80000000;
defparam prom_inst_13.INIT_RAM_0A = 256'hF0003FF83F87807F80007C00007FFFFFE00000007FFFFFF1C01001FFBE51AFFF;
defparam prom_inst_13.INIT_RAM_0B = 256'h1F03F000FFF81F87C07E000FFF03F83F0FC000FFF07F83E0FF0003FF87F03F0F;
defparam prom_inst_13.INIT_RAM_0C = 256'hFFFC8000024800007FFFFFE0007FFF00000FFFFE007FF81FC0F8DF001FFF83FC;
defparam prom_inst_13.INIT_RAM_0D = 256'h0000000FFFFFF90000000000FFFFFFBC000000004F3FFFA412F52060000003FF;
defparam prom_inst_13.INIT_RAM_0E = 256'h000007FFFFF21FB0000003FFFFFD0000000000FFFFFE40000000003FFFFFFE00;
defparam prom_inst_13.INIT_RAM_0F = 256'h000003FFFFFFFFF0000003FFFFFFFFF8000003FFFFFFFFF8000003FFFFFF7FF0;
defparam prom_inst_13.INIT_RAM_10 = 256'h000FFFFFFFFFFC000000FFFFFFFFFF0000001FFFFFFFFFE0000007FFFFF6FFF8;
defparam prom_inst_13.INIT_RAM_11 = 256'hF000FFFF0000007FFFFC00FFFF0000007FFFFC00FFFC000001FFFFF817FFC000;
defparam prom_inst_13.INIT_RAM_12 = 256'hFFFFF0000FFFF8000001FFFFFF000FFFF8000001FFFFFF0003FFF0000007FFFF;
defparam prom_inst_13.INIT_RAM_13 = 256'hFFFFF800001FFFE000003FFFFFC00003FFFE000001FFFFFF00007FFFC000000F;
defparam prom_inst_13.INIT_RAM_14 = 256'hFFFFE000007FFFC000007FFFFC000007FFFC000007FFFFF000001FFFF800001F;
defparam prom_inst_13.INIT_RAM_15 = 256'h7FFFFF803FFFFF80000003FFFFE000FFFFFF0000003FFFFE00006FFFFC000003;
defparam prom_inst_13.INIT_RAM_16 = 256'h007FFFFFFFFF800000000007FFFFFFFFFFF0000000007FFFFFFFFFFE00000000;
defparam prom_inst_13.INIT_RAM_17 = 256'hACCE6A644A492AD96B76924EA54A54CCC997291B13B2A488D908001000000000;
defparam prom_inst_13.INIT_RAM_18 = 256'hD448A6766664C95996ECD991A454D9899999A52D5936A5492AA44C8C936A6CC4;
defparam prom_inst_13.INIT_RAM_19 = 256'hCCCECCCC0A4ADD4C4AD7B672A4288DCCCC999966664ECC446E6766733B337666;
defparam prom_inst_13.INIT_RAM_1A = 256'h07F3FFFFFC00400FF7FFFFE000200FFFFFFFE000003FFFFFFB320000009FFFDD;
defparam prom_inst_13.INIT_RAM_1B = 256'hEFFF000003FFFF27FFC00603FBFF81FF803F07F1FF07FF007F07E1FFFFFF003E;
defparam prom_inst_13.INIT_RAM_1C = 256'h000000007FFFFFFFF000000003FFFFFFF800000001FFFFFF80000000003FFFFF;
defparam prom_inst_13.INIT_RAM_1D = 256'h21FFFFFF000000000FFFFFFFF00000000003FFFFFFFFFB000000001FFFFFFFFF;
defparam prom_inst_13.INIT_RAM_1E = 256'h0000014F8D90000000001E948007E36400000002000006DFFFFC000000000000;
defparam prom_inst_13.INIT_RAM_1F = 256'h000020218482000000000000013002000000000010FB5F6C0000000965FDC800;
defparam prom_inst_13.INIT_RAM_20 = 256'h8001DFFA1002D210ABFE8063520008D4FFFC000400000200001FFD0000001000;
defparam prom_inst_13.INIT_RAM_21 = 256'h07E3FFFFF401FC1F99FFFE007807FFFFFC0000001FFFFFFFF180000FFFF000FE;
defparam prom_inst_13.INIT_RAM_22 = 256'hFFFFC03F807C7FFFFFE00FC07E7FFFFFC03FE0F87FEFFF801F03F8FFFFFF00FF;
defparam prom_inst_13.INIT_RAM_23 = 256'h1FE7FFFFFF003301FE7FFFFFF006703FCFFCFFFE00FE0FF1FFFFFFC07F00FCFF;
defparam prom_inst_13.INIT_RAM_24 = 256'hDC0FF1FFFFFFF003303FE7FFFFFF8008C0FF9FFFFFFE003703FCFFFFFFE00030;
defparam prom_inst_13.INIT_RAM_25 = 256'h701FEFFFE3FFFC01BC07F3FFF1FFFC00FE07F9FFFDFFFE00FE07F1FFEFFFF801;
defparam prom_inst_13.INIT_RAM_26 = 256'hFBFFC01FFFE00FC07F9FFC00FFFE00FE07F9FF801FFFC00BC0FF3FF803FFF003;
defparam prom_inst_13.INIT_RAM_27 = 256'h1FFF800001FFFFF8003FFF800001FFFFF8007FFF800401FFFFF001FFFC00F80F;
defparam prom_inst_13.INIT_RAM_28 = 256'hFFFF8003FFE000003FFFFFF80007FFC00001FFFFFFC0003FFC00000FFFFFF000;
defparam prom_inst_13.INIT_RAM_29 = 256'hFFFF0000005FFC00001FFFFFEA0000009EC000007FFFFFFA8000FFF800001FFF;
defparam prom_inst_13.INIT_RAM_2A = 256'hFFFFF00003FFF800007FFFFFFF80000FFFC00003FFFFFFF8000077FE00001FFF;
defparam prom_inst_13.INIT_RAM_2B = 256'hFE000800001FFF80003FFFFF8EC00003FFF80001FFFFFFFC00001FFF80000FFF;
defparam prom_inst_13.INIT_RAM_2C = 256'h001FFE0001FFF00007FFFE0007FE0001FFF00007F7FE0007F80007FFF0001FFF;
defparam prom_inst_13.INIT_RAM_2D = 256'hFF000FFE0000FFFFF80003FF0007FF80001FFFFFE0001FFC0007FF80007FFFFC;
defparam prom_inst_13.INIT_RAM_2E = 256'h000003FFFFFFE0001FFE000FF80000FFFFFF00007FA003FE00007FFFFFF0000F;
defparam prom_inst_13.INIT_RAM_2F = 256'h000000002FFFFFFFFFFFFD000000007FFFF800BFFF8000000003FFFFFFF00000;
defparam prom_inst_13.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000001E79E10;
defparam prom_inst_13.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_13.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_13.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_13.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_13.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_13.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_13.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_13.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_13.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_13.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_13.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_13.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_13.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_13.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_13.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

pROM prom_inst_14 (
    .DO({prom_inst_14_dout_w[30:0],prom_inst_14_dout[7]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_14.READ_MODE = 1'b0;
defparam prom_inst_14.BIT_WIDTH = 1;
defparam prom_inst_14.RESET_MODE = "SYNC";
defparam prom_inst_14.INIT_RAM_00 = 256'h0000000000000000000000000000000000000000000000000000000000005547;
defparam prom_inst_14.INIT_RAM_01 = 256'h000000000000000000000000019290281E929010A03A4A406280E929010A0384;
defparam prom_inst_14.INIT_RAM_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_20 = 256'h07F80007FFFBFFFC07F00001FFFFFFFC1FE00000007FFE07FFC00F804FE8003F;
defparam prom_inst_14.INIT_RAM_21 = 256'hFC3FFC0001FFF1FFE07FE0001FFFFFFF81FF80007FFFFFFF01FE0000FFFFFFFC;
defparam prom_inst_14.INIT_RAM_22 = 256'hFFFFFFFFFE0001FFFFFFFFFFC0003FFF7FFFFFF80003FFFFFFFFFF80001FFEFF;
defparam prom_inst_14.INIT_RAM_23 = 256'h000007FFF57FFFE00000FFFFCFFFF800003FFFFFFFFF00000FFFFFFFFFE00007;
defparam prom_inst_14.INIT_RAM_24 = 256'hFF00000001FFFFFFFE00000000FFFFFFF80000003FFFFFFFE000001FFFFFFFFF;
defparam prom_inst_14.INIT_RAM_25 = 256'hF00000000FFFFFFFFC00000001FFFFFFFF00000000FFFFFFFF00000001FFFFFF;
defparam prom_inst_14.INIT_RAM_26 = 256'h000003FFFFFFFFE00000000FFFFFFFFC00000003FFFFFFFFC00000003FFFFFFF;
defparam prom_inst_14.INIT_RAM_27 = 256'hAFFFFFFFA0000000F7FFFFFFFF80000000AFFFFFFFFF800000005FFFFFFFFE00;
defparam prom_inst_14.INIT_RAM_28 = 256'hE0000022FFFFFFFFFFE0000016FDFFFFFFFFC00000056AAFFFFFFFF000000028;
defparam prom_inst_14.INIT_RAM_29 = 256'h00FFF801FFFFFC00002FFFDAFFFFFF8000017FFFF7FFFFFC00000CFD7FFFFFFF;
defparam prom_inst_14.INIT_RAM_2A = 256'hF8001FFFFE000007FFC003FFFFF000007FF8003FFFFE00000FFF800FFFFFC000;
defparam prom_inst_14.INIT_RAM_2B = 256'hFFF000003FFFC001FFFFF000003FFF8001FFFFF000007FFE0003FFFFC00001FF;
defparam prom_inst_14.INIT_RAM_2C = 256'h80001FFFFFE00003FFFC4000FFFFFC00003FFFFE000FFFFF800003FFFFD001FF;
defparam prom_inst_14.INIT_RAM_2D = 256'h07FFF800001FFFFFC00003FFF000007FFFFF00001FFFE00001FFFFFC00003FFF;
defparam prom_inst_14.INIT_RAM_2E = 256'hE00003FFF00000FFFFFFC00007FFF00001FFFFFF800007FFF00003FFFFFFC000;
defparam prom_inst_14.INIT_RAM_2F = 256'hFFFF800007FFF00003FFFFFFC00003FFF80000FFFFFFE00003FFF80000FFFFFF;
defparam prom_inst_14.INIT_RAM_30 = 256'h0FFFFFFFC00003FFE00003FFFFFF800007FFC00003FFFFFF800007FFE00003FF;
defparam prom_inst_14.INIT_RAM_31 = 256'h00000BFFFFFFF000007FE00007FFFFFFE00001FF800007FFFFFFC00003FF8000;
defparam prom_inst_14.INIT_RAM_32 = 256'h000000001FFFFFFFFE00000000000FFFFFFFFC000000000007FFFFFFF800001B;
defparam prom_inst_14.INIT_RAM_33 = 256'hFFFF5000000002FFFFFFFFFF0000000003FFFFFFFFE80000000001FFFFFFFF00;
defparam prom_inst_14.INIT_RAM_34 = 256'h000A00FFFFF000007F800FFFFFFE000003FFFFEB01FFFFFE4400000007FFFFFF;
defparam prom_inst_14.INIT_RAM_35 = 256'hFFE000005E00000FFFFFF000001FFFF0007FFFFF00000001FFFFFFFFC00007FF;
defparam prom_inst_14.INIT_RAM_36 = 256'h007FFFFFFFE00000000007FFFFFFFF00000000000FFFFFFFE00000000003FFFF;
defparam prom_inst_14.INIT_RAM_37 = 256'h0001FFFFFFFFFFFF80000003FFFFFFFFFFFE0000001FFF7FFFFFFFFE00000000;
defparam prom_inst_14.INIT_RAM_38 = 256'hF0000000065FFFFFFFFFE000000000BFFFFFFFFFC00000007FFFFFFFFFFF8000;
defparam prom_inst_14.INIT_RAM_39 = 256'h3FFF000000000487FFFFFFFFF800000008C17FFFFFFFF80000000003FFFFFFFF;
defparam prom_inst_14.INIT_RAM_3A = 256'h0000001FFFFC1FFFF000000EFFFFE3FFFE0000007FFFFFFFFFE0000001FFFFF0;
defparam prom_inst_14.INIT_RAM_3B = 256'h07FFFFFFFFFF00000007FFFFFFFFFC00000007FFFFFFFFE00000007FFFE1FFFE;
defparam prom_inst_14.INIT_RAM_3C = 256'hFFE00000000FFFFFFFFFC00000003FFFFFFFFFFE00000003FFFFFFFFFF000000;
defparam prom_inst_14.INIT_RAM_3D = 256'h001FFFFFFFFF00000000FFFFFFFFFF00000001FFFFFFFFFFC0000000FFFFFFFF;
defparam prom_inst_14.INIT_RAM_3E = 256'hFFFFFFF8000003FFFFFFFFFF0000003FFFFFFFFFF8000007FFFFFFFFFFE00000;
defparam prom_inst_14.INIT_RAM_3F = 256'hE01FFF00007FFFFFE03FFF800007FFFFF03FFF8000107FFFFFFFFFE00001FFFF;

pROM prom_inst_15 (
    .DO({prom_inst_15_dout_w[30:0],prom_inst_15_dout[7]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_15.READ_MODE = 1'b0;
defparam prom_inst_15.BIT_WIDTH = 1;
defparam prom_inst_15.RESET_MODE = "SYNC";
defparam prom_inst_15.INIT_RAM_00 = 256'hF001FF0000FF9FFFF003FF80007F9FFFF003FF0000FFFFFFF00FFF00007FFFFF;
defparam prom_inst_15.INIT_RAM_01 = 256'h01FE00063FFF83FE001FE0003FFFFC7FC007FC0001FFFF1FE003FF0001FFFF3F;
defparam prom_inst_15.INIT_RAM_02 = 256'h3F87FFF03FC00FF0007F07FFF03F9F0FF000003FFFE0FFFC3FC000E07FFC1FE1;
defparam prom_inst_15.INIT_RAM_03 = 256'h7F8000FF9F87FFC0FFF83F0001FFFF3FFE07FFC1F8000FFF7FFFC0FFF83FC000;
defparam prom_inst_15.INIT_RAM_04 = 256'hFF8FC0007FFF381F1F07FFC1F8000FFF9F81CFE0FFF87E0000FF87C1FFF03FF8;
defparam prom_inst_15.INIT_RAM_05 = 256'hFFF80001FFFFF0F0F038FFFC7C0001FFFFFE0187C3FFF1F8000FFFFF0F80FC1F;
defparam prom_inst_15.INIT_RAM_06 = 256'hF800007FFFF83FF81FFFFFF00003FFFFE0FC001FFFFFF000007FFFFC30F019FF;
defparam prom_inst_15.INIT_RAM_07 = 256'hF000001FFFFFFFFFFFFFFE000003FFFFFEFFFFFFFFF800001FFFFF1FBF0FFFFF;
defparam prom_inst_15.INIT_RAM_08 = 256'hFFC000000000D3FFFFFFFFF00000001FFFFFFFFFFFFC0000003FFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_09 = 256'h011FFFCFFC00001FFFFFFFFFFE0000000003FFFFFFFFFF80000000007FFFFFFF;
defparam prom_inst_15.INIT_RAM_0A = 256'h0FFFC007FFF800007FFF83FFFF8000001FFFFFFF8000000E3FEFFE0041AE5000;
defparam prom_inst_15.INIT_RAM_0B = 256'hE0000FFF0007FFF80001FFF000FFFFC0003FFF000FFFFC0000FFFC007FFFC000;
defparam prom_inst_15.INIT_RAM_0C = 256'h00037FFFFDB7FFFF8000001FFF8000FFFFF00001FF8007FFFF0000FFE0007FFF;
defparam prom_inst_15.INIT_RAM_0D = 256'hFFFFFFF0000006FFFFFFFFFF00000043FFFFFFFFB0C0005BED0ADF9FFFFFFC00;
defparam prom_inst_15.INIT_RAM_0E = 256'hFFFFF800000DE04FFFFFFC000002FFFFFFFFFF000001BFFFFFFFFFC0000001FF;
defparam prom_inst_15.INIT_RAM_0F = 256'hFFFFFC000000000FFFFFFC0000000007FFFFFC0000000007FFFFFC000000800F;
defparam prom_inst_15.INIT_RAM_10 = 256'hFFF00000000003FFFFFF0000000000FFFFFFE0000000001FFFFFF80000090007;
defparam prom_inst_15.INIT_RAM_11 = 256'h0FFF0000FFFFFF800003FF0000FFFFFF800003FF0003FFFFFE000007E8003FFF;
defparam prom_inst_15.INIT_RAM_12 = 256'h00000FFFF00007FFFFFE000000FFF00007FFFFFE000000FFFC000FFFFFF80000;
defparam prom_inst_15.INIT_RAM_13 = 256'h000007FFFFE0001FFFFFC000003FFFFC0001FFFFFE000000FFFF80003FFFFFF0;
defparam prom_inst_15.INIT_RAM_14 = 256'h00001FFFFF80003FFFFF800003FFFFF80003FFFFF800000FFFFFE00007FFFFE0;
defparam prom_inst_15.INIT_RAM_15 = 256'h8000007FC000007FFFFFFC00001FFF000000FFFFFFC00001FFFF900003FFFFFC;
defparam prom_inst_15.INIT_RAM_16 = 256'hFF80000000007FFFFFFFFFF800000000000FFFFFFFFF800000000001FFFFFFFF;
defparam prom_inst_15.INIT_RAM_17 = 256'h5331959BB5B6D52694896DB15AB5AB333668D6E4EC4D5B7726F7001FFFFFFFFF;
defparam prom_inst_15.INIT_RAM_18 = 256'h2BB75989999B36A66913266E5BAB267666665AD2A6C95AB6D55BB3736C95933B;
defparam prom_inst_15.INIT_RAM_19 = 256'h33313333F5B522B3B528498D5BD772333366669999B133BB9198998CC4CC8999;
defparam prom_inst_15.INIT_RAM_1A = 256'hF800000003FFFFF00000001FFFFFF00000001FFFFFC0000004CDFFFFFF600022;
defparam prom_inst_15.INIT_RAM_1B = 256'h1000FFFFFC0000D8003FFFFC00007E007FFFF80000F800FFFFF800000000FFFF;
defparam prom_inst_15.INIT_RAM_1C = 256'hFFFFFFFF800000000FFFFFFFFC00000007FFFFFFFE0000007FFFFFFFFFC00000;
defparam prom_inst_15.INIT_RAM_1D = 256'hDE000000FFFFFFFFF00000000FFFFFFFFFFC0000000004FFFFFFFFE000000000;
defparam prom_inst_15.INIT_RAM_1E = 256'hFFFFFEB0726FFFFFFFFFE16B7FF81C9BFFFFFFFDFFFFF9200003FFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_1F = 256'hFFFFDFDE7B7DFFFFFFFFFFFFFECFFDFFFFFFFFFFEF04A093FFFFFFF69A0237FF;
defparam prom_inst_15.INIT_RAM_20 = 256'h7FFE2005EFFD2DEF54017F9CADFFF72B0003FFFBFFFFFDFFFFE002FFFFFFEFFF;
defparam prom_inst_15.INIT_RAM_21 = 256'hF80000000BFFFFE0000001FFFFF8000003FFFFFFE00000000E7FFFF0000FFF01;
defparam prom_inst_15.INIT_RAM_22 = 256'h00003FFFFF800000001FFFFF800000003FFFFF000010007FFFFC00000000FFFF;
defparam prom_inst_15.INIT_RAM_23 = 256'hE000000000FFFFFE000000000FFFFFC000030001FFFFF0000000003FFFFF0000;
defparam prom_inst_15.INIT_RAM_24 = 256'hFFF0000000000FFFFFC0000000007FFFFF0000000001FFFFFC000000001FFFFF;
defparam prom_inst_15.INIT_RAM_25 = 256'hFFE000001C0003FFFFF800000E0003FFFFF80000020001FFFFF80000100007FF;
defparam prom_inst_15.INIT_RAM_26 = 256'h00003FE0001FFFFF800003FF0001FFFFF800007FE0003FFFFF000007FC000FFF;
defparam prom_inst_15.INIT_RAM_27 = 256'hE0007FFFFE000007FFC0007FFFFE000007FF80007FFFFE00000FFE0003FFFFF0;
defparam prom_inst_15.INIT_RAM_28 = 256'h00007FFC001FFFFFC0000007FFF8003FFFFE0000003FFFC003FFFFF000000FFF;
defparam prom_inst_15.INIT_RAM_29 = 256'h0000FFFFFFA003FFFFE0000015FFFFFF613FFFFF800000057FFF0007FFFFE000;
defparam prom_inst_15.INIT_RAM_2A = 256'h00000FFFFC0007FFFF800000007FFFF0003FFFFC00000007FFFF8801FFFFE000;
defparam prom_inst_15.INIT_RAM_2B = 256'h01FFF7FFFFE0007FFFC00000713FFFFC0007FFFE00000003FFFFE0007FFFF000;
defparam prom_inst_15.INIT_RAM_2C = 256'hFFE001FFFE000FFFF80001FFF801FFFE000FFFF80001FFF807FFF8000FFFE000;
defparam prom_inst_15.INIT_RAM_2D = 256'h00FFF001FFFF000007FFFC00FFF8007FFFE000001FFFE003FFF8007FFF800003;
defparam prom_inst_15.INIT_RAM_2E = 256'hFFFFFC0000001FFFE001FFF007FFFF000000FFFF805FFC01FFFF8000000FFFF0;
defparam prom_inst_15.INIT_RAM_2F = 256'hFFFFFFFFD0000000000002FFFFFFFF800007FF40007FFFFFFFFC0000000FFFFF;
defparam prom_inst_15.INIT_RAM_30 = 256'h00000000000000000000000000000000000000000000000000000000011861EF;
defparam prom_inst_15.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_15.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce)
);
MUX2 mux_inst_0 (
  .O(dout[0]),
  .I0(prom_inst_0_dout[0]),
  .I1(prom_inst_1_dout[0]),
  .S0(dff_q_0)
);
MUX2 mux_inst_1 (
  .O(dout[1]),
  .I0(prom_inst_2_dout[1]),
  .I1(prom_inst_3_dout[1]),
  .S0(dff_q_0)
);
MUX2 mux_inst_2 (
  .O(dout[2]),
  .I0(prom_inst_4_dout[2]),
  .I1(prom_inst_5_dout[2]),
  .S0(dff_q_0)
);
MUX2 mux_inst_3 (
  .O(dout[3]),
  .I0(prom_inst_6_dout[3]),
  .I1(prom_inst_7_dout[3]),
  .S0(dff_q_0)
);
MUX2 mux_inst_4 (
  .O(dout[4]),
  .I0(prom_inst_8_dout[4]),
  .I1(prom_inst_9_dout[4]),
  .S0(dff_q_0)
);
MUX2 mux_inst_5 (
  .O(dout[5]),
  .I0(prom_inst_10_dout[5]),
  .I1(prom_inst_11_dout[5]),
  .S0(dff_q_0)
);
MUX2 mux_inst_6 (
  .O(dout[6]),
  .I0(prom_inst_12_dout[6]),
  .I1(prom_inst_13_dout[6]),
  .S0(dff_q_0)
);
MUX2 mux_inst_7 (
  .O(dout[7]),
  .I0(prom_inst_14_dout[7]),
  .I1(prom_inst_15_dout[7]),
  .S0(dff_q_0)
);
endmodule //GSrom_test
