//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.10.03 (64-bit)
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Mon Dec  9 21:37:33 2024

module rom_gs105b (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [14:0] ad;

wire lut_f_0;
wire lut_f_1;
wire [30:0] prom_inst_0_dout_w;
wire [0:0] prom_inst_0_dout;
wire [30:0] prom_inst_1_dout_w;
wire [0:0] prom_inst_1_dout;
wire [30:0] prom_inst_2_dout_w;
wire [1:1] prom_inst_2_dout;
wire [30:0] prom_inst_3_dout_w;
wire [1:1] prom_inst_3_dout;
wire [30:0] prom_inst_4_dout_w;
wire [2:2] prom_inst_4_dout;
wire [30:0] prom_inst_5_dout_w;
wire [2:2] prom_inst_5_dout;
wire [30:0] prom_inst_6_dout_w;
wire [3:3] prom_inst_6_dout;
wire [30:0] prom_inst_7_dout_w;
wire [3:3] prom_inst_7_dout;
wire [30:0] prom_inst_8_dout_w;
wire [4:4] prom_inst_8_dout;
wire [30:0] prom_inst_9_dout_w;
wire [4:4] prom_inst_9_dout;
wire [30:0] prom_inst_10_dout_w;
wire [5:5] prom_inst_10_dout;
wire [30:0] prom_inst_11_dout_w;
wire [5:5] prom_inst_11_dout;
wire [30:0] prom_inst_12_dout_w;
wire [6:6] prom_inst_12_dout;
wire [30:0] prom_inst_13_dout_w;
wire [6:6] prom_inst_13_dout;
wire [30:0] prom_inst_14_dout_w;
wire [7:7] prom_inst_14_dout;
wire [30:0] prom_inst_15_dout_w;
wire [7:7] prom_inst_15_dout;
wire dff_q_0;

LUT2 lut_inst_0 (
  .F(lut_f_0),
  .I0(ce),
  .I1(ad[14])
);
defparam lut_inst_0.INIT = 4'h2;
LUT2 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(ad[14])
);
defparam lut_inst_1.INIT = 4'h8;
pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[30:0],prom_inst_0_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 1;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hFFFFFFFFFFCC206EB424D628274C536CFCD757FFFFFFDDC00EF9FFFFFFFFFF3B;
defparam prom_inst_0.INIT_RAM_01 = 256'h86590A318601111F8F742E55E7D175365334FFFF8509FF00093A6AF06BC60E2B;
defparam prom_inst_0.INIT_RAM_02 = 256'hFFFFFFFFFFFEABA49C2B671A40657EAAD1414E5BC7744FF32002A50A94C4EEEE;
defparam prom_inst_0.INIT_RAM_03 = 256'h4BE967E0203D2101E9E03D3B4EEF3BB6524933A7AA9A1469A0006BEB105EBABB;
defparam prom_inst_0.INIT_RAM_04 = 256'h4EAE89420484E2A3A48B4AA2939102499F8B4A5C9725C9D2E424B97E90917E9E;
defparam prom_inst_0.INIT_RAM_05 = 256'h4E73A828282821CFF48AFEFFBFD39C931498DC8BFFFFCFB9FE974FB4E7FA7464;
defparam prom_inst_0.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFF2AE7D391439C22039CE7C1F14C27D3CF8B4C9F4FA5E949C9F;
defparam prom_inst_0.INIT_RAM_07 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_0.INIT_RAM_08 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_0.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF52C3BF2EEA5976A0;
defparam prom_inst_0.INIT_RAM_0A = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_0.INIT_RAM_0B = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_0.INIT_RAM_0C = 256'h8AAA8ACAA984D1AB4A476E302B218158714933894605648039C4808508B72550;
defparam prom_inst_0.INIT_RAM_0D = 256'hD74E6EB4D374524F7C67995AF1B5AAD8A9290EECC450A488015200429CEA8A8A;
defparam prom_inst_0.INIT_RAM_0E = 256'h42F9DA273F39F5CFADDB5D39B2FD67D7EB3ED24A5A5DB5D39BD7DDB4E6AE7B76;
defparam prom_inst_0.INIT_RAM_0F = 256'h511AA834B0237051DC342AD0556ECFF1D718F58BA4D53169A36AC7558A20A022;
defparam prom_inst_0.INIT_RAM_10 = 256'h756BE6BA793FAC098212934DFCDD2AA5475D26725D0D87DD9A2E60D5D91C3C31;
defparam prom_inst_0.INIT_RAM_11 = 256'hF679A4D008321E649E6CC2185E6F19A6CD972A1164AB7AEBB11ABADAAA69E59A;
defparam prom_inst_0.INIT_RAM_12 = 256'hEE5E3CEAE447ACF4999E03DFC3FB2AB35206853A2DEF7AD6EDEF5147AD687F69;
defparam prom_inst_0.INIT_RAM_13 = 256'h32AA03F1316218DA877B003AF60075F700EBEE01D76C03AE6E075C370EB800D1;
defparam prom_inst_0.INIT_RAM_14 = 256'h16126C14A6015FC4C5886305553FFC4C58901FC4C588418AAAAAAAAA7B58B06D;
defparam prom_inst_0.INIT_RAM_15 = 256'h7CCC87D1CD367DF697C26E9AF66E2EA2D24D228AD07BEFAD97B5DBC540475F13;
defparam prom_inst_0.INIT_RAM_16 = 256'hFFFFFFD1AA2D000000800E03830C4C169325C112DA4452B35B86B20BFCF4E945;
defparam prom_inst_0.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_0.INIT_RAM_18 = 256'h0828005F5DD7D55F75F7F60A082880357FD74A888F7FCA0D70BC8A8877D5F5D6;
defparam prom_inst_0.INIT_RAM_19 = 256'h02757D7D7D7F57F55FFF5555555FFD57F5F5F7DC22222228A0A02AAAAA0A0822;
defparam prom_inst_0.INIT_RAM_1A = 256'h015B1D1650346E59F1ADD04F7224F63030EBD99BCBA495531658160002741600;
defparam prom_inst_0.INIT_RAM_1B = 256'h65EF332A96773F49F3CDD34F0B199C9376E9F673A8FA2552A9441D9A4CC6AD97;
defparam prom_inst_0.INIT_RAM_1C = 256'h3A7FC88FC6BEBAE7E7F83DEC3D5CBD55FE7349A74D3DF724E92EE943CB2E8EA9;
defparam prom_inst_0.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF38E7CFBAE9C1;
defparam prom_inst_0.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_0.INIT_RAM_20 = 256'h453F1CF29FF6C20E1FB611C3F6C839FB6473F6C8502D97827565000B1113BBAB;
defparam prom_inst_0.INIT_RAM_21 = 256'hF30C77A6FD77E9BF4DFA6FFEEDFB4F37075B6414FC73C29FF6C8A7E0E794FFB6;
defparam prom_inst_0.INIT_RAM_22 = 256'hE66648857332257D5757BAACBDD57AAAB21FF99AF8E88EA47559FA32D1DD643F;
defparam prom_inst_0.INIT_RAM_23 = 256'hBAA54822BAA442BE9BE9D2DD2EC9D044AEC94457D3B5BAB20B644AEC82257C76;
defparam prom_inst_0.INIT_RAM_24 = 256'hAC9918457D3B5BAD45714CCAC95A88C232576978EF8E46654CACC5723B232574;
defparam prom_inst_0.INIT_RAM_25 = 256'h8B122C82C48B146399D2F55B2B657115AA99590AFA6FA74B7697B59B32B8AC95;
defparam prom_inst_0.INIT_RAM_26 = 256'hCB632D16B2C5ACB630B16B2C518E6B6D46DAEA2C8B162D122D8B160B162C8B44;
defparam prom_inst_0.INIT_RAM_27 = 256'hFEF65556A32C959D6E8AB21FF986E7031B69E30B2B2C48CB448CB2B2C48C2C48;
defparam prom_inst_0.INIT_RAM_28 = 256'hD1E2D10AA858A45885B6A9445885162C162C42DD9558ECB3F5557BAAC87FE61B;
defparam prom_inst_0.INIT_RAM_29 = 256'h88536D518B8B10B246582465885B52E8B10AA1162058A16C616285922C48B442;
defparam prom_inst_0.INIT_RAM_2A = 256'h5D5AD4BB8658859030B14B2C50B51962055432C52CB442D2AB2D10AA46589185;
defparam prom_inst_0.INIT_RAM_2B = 256'h554E8B458B10BF162174A2C42F41621756C59E8B122C50BD16205D22C42F4588;
defparam prom_inst_0.INIT_RAM_2C = 256'h478B122D10AD16085562C50AF1620555A96BA2C582C42BD1621558B442BC5821;
defparam prom_inst_0.INIT_RAM_2D = 256'h14EB2C42CB185885BAE2C42C8DB16F2E2C52CB142F865881742CB10BC1962175;
defparam prom_inst_0.INIT_RAM_2E = 256'h285A8CB1028ADE969C32C50C2C42B971621550CB442B965821554F51960B1962;
defparam prom_inst_0.INIT_RAM_2F = 256'hFD23A805278A10FD823AC452FB57FF28AD74EE879C6589596885A8CB042C9596;
defparam prom_inst_0.INIT_RAM_30 = 256'h38EFFDEF3FEFFFFFF9FE7FDFE7F08A8053440C7EC0540205CFFBFFFDFE9FF7F9;
defparam prom_inst_0.INIT_RAM_31 = 256'h3F67F95FFFFFFFDFEFFFFFFFFFE0CEB1431FB07FD7114B3A840C7EE5FEFBD7FF;
defparam prom_inst_0.INIT_RAM_32 = 256'h1061765C120EB8A38BA039F3BFFFFFFFFFFFFFFFFFFFC0A840C7EC6888C56284;
defparam prom_inst_0.INIT_RAM_33 = 256'hF7F9FF7FFF823AC51100299D4200801FEFF5DCFFBFCFFBFBFD3FEFF3FEFE09D6;
defparam prom_inst_0.INIT_RAM_34 = 256'hF9FDFE9FF7F9FF7F9FC13AC51431FB029075082043F722B8EE7FDFE7F6FFFE9F;
defparam prom_inst_0.INIT_RAM_35 = 256'h4FFFEFF7FC11D420810FD80299D628A18A1FB94FFBFCFFBFCFFFEB39FF7F9FF7;
defparam prom_inst_0.INIT_RAM_36 = 256'h7F7FB7F00EB1450C50FDC9003AC5143143F729FF7F9FF7F9FDAE3B9FF7F9FF7F;
defparam prom_inst_0.INIT_RAM_37 = 256'h823A84102163F712B6758A286287EE253FEFF3FEFF3FEFFFEBB9FF7F9FF7F9FF;
defparam prom_inst_0.INIT_RAM_38 = 256'hA1FB89202758A286287EE253FEFF3FEFF3FEFE679DCFFBFCFFBFCFEDFFFDFEFF;
defparam prom_inst_0.INIT_RAM_39 = 256'h510C50FDC4A7FDFE7FDFE7FDFE7FFF31CFFBFCFFBFCFFBFCFEFF4FE49D628A18;
defparam prom_inst_0.INIT_RAM_3A = 256'h7FDFE7FDFE7FFB0EE7FDFE7FDFE7FDFD3FFFBFDFF82750820042C7EE24E8EB14;
defparam prom_inst_0.INIT_RAM_3B = 256'hFF7F9FF7F9FF7F9FF7F7FB7F68EB14510C50FDC49023AC51443143F711A7FDFE;
defparam prom_inst_0.INIT_RAM_3C = 256'hEFF003A8410020163F71232758A28862287EE253FEFF3FEFF3FEFF3FEFFFE2B9;
defparam prom_inst_0.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFFBFCFFBFCFFBFCFEDFFFDF;
defparam prom_inst_0.INIT_RAM_3E = 256'h6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6;
defparam prom_inst_0.INIT_RAM_3F = 256'hDB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6DB6D;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[30:0],prom_inst_1_dout[0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 1;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h40240240244F03A40094CFD67EA7C0B0559BCCFDDD801541027FFF84FFFF0903;
defparam prom_inst_1.INIT_RAM_01 = 256'hD252D8E8A8FA2A3A8A8EB3A266A2BB3332A219EA2BB3332A61C3E2589A402402;
defparam prom_inst_1.INIT_RAM_02 = 256'h1F17DE63FD814FEF3FED28360801DF4211DA4B6AAC93B928AA8A8AA8CA8D62B0;
defparam prom_inst_1.INIT_RAM_03 = 256'h6866E00451A57146FB1810027715A540A7751810027713321A0375332180371F;
defparam prom_inst_1.INIT_RAM_04 = 256'h990F01BEADD4223D1B8BF71F1888F31533219A711349A69D86800A3C0088A98B;
defparam prom_inst_1.INIT_RAM_05 = 256'h96DBC23D1F5FAE8B3A3B2A33F98DDDF98F75C89DFC0EF401EFA498012925FFE9;
defparam prom_inst_1.INIT_RAM_06 = 256'hFE2F73F8FDEFE2C2F4775FAEF83D1D9990C01B88DC7E8DE28E3E02057E2DB79F;
defparam prom_inst_1.INIT_RAM_07 = 256'h5D31D76BFFC98531004004FE39F4744555A37BEDCF6DFDFC5BEDEFE3F7BF8BDC;
defparam prom_inst_1.INIT_RAM_08 = 256'h1F7AF57F7E4EEB71F0493F527BF3FAB51ACCF846AB51ACCF846AFBEBE06FC3D4;
defparam prom_inst_1.INIT_RAM_09 = 256'hE27D78276D3FAD319BFAFD763B913FDFC427EBB5F268FFFF4D3F1102BC799930;
defparam prom_inst_1.INIT_RAM_0A = 256'hFEDA66E9EB7B4D38A13849FC93E93D8AD24D3E5154450CB831B0CFDEE98C2642;
defparam prom_inst_1.INIT_RAM_0B = 256'h7E7F462F99AAA8A8ECECFAEBDDCD34E5F35FC9B69CFFB699BA7ADED276C90793;
defparam prom_inst_1.INIT_RAM_0C = 256'h81F6BD37DBBE3D39BAB595B34FD9A3F0BD0479E08F3C7B2392BEAAF928A5EBAE;
defparam prom_inst_1.INIT_RAM_0D = 256'h042615B1AEF2EC6A3DBDB1ADF5A151EDE1CDF6ECCFBA7FDD1FB7E823CF047A89;
defparam prom_inst_1.INIT_RAM_0E = 256'h7AD7646A338828A068AAB43E77322981602885A1154551A05E86BCF3CF38E38E;
defparam prom_inst_1.INIT_RAM_0F = 256'h9477652492492492FDBF6EEBFF7EFDFBEFBEFAFDF5FBF7A8AA0D769E31EFB6CC;
defparam prom_inst_1.INIT_RAM_10 = 256'hDD13AFCC78F5C460C74EC576ECCEBBD6F8F7ED26ECCEBBD6F8EE6749D7C778E7;
defparam prom_inst_1.INIT_RAM_11 = 256'h91644A611A519EE49FEE1BA7C72AEA322EDBE0E3D48B225308D28CFE8ABD7EBA;
defparam prom_inst_1.INIT_RAM_12 = 256'hCD8072D85BCCCCF031BB333DF0890F0ED0BBFEE1319029DB9D594645DB1C1C1A;
defparam prom_inst_1.INIT_RAM_13 = 256'h1A01E50350224F8AF9E667CE7FDBAFCB9CDEE7F962E7A7FF2E737BAFD57DA96A;
defparam prom_inst_1.INIT_RAM_14 = 256'h1D78D46D683B6A47EECF3D8DBE318C13140F2D1D1BEEAA8201A81081CD021029;
defparam prom_inst_1.INIT_RAM_15 = 256'hBD60000DDBD787D5976DAB0704561105677CFF111FF3FF7518DD5DA7618E3DC9;
defparam prom_inst_1.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF555A54352A805DD8B5E;
defparam prom_inst_1.INIT_RAM_17 = 256'h0000FFFFFFFFFFFFFFFF0000FFFFFFFFFFFFF3F8FFFFFE181897FFFA569392D4;
defparam prom_inst_1.INIT_RAM_18 = 256'h00000000000000000000FFFFFFFFFFFF000000000001038041C1FC0000000000;
defparam prom_inst_1.INIT_RAM_19 = 256'h00000113AAAABBB0FBFFFFFFFB2FAEC3FFFFFFFFFFCFAB02FFFFFFFF346AAAAA;
defparam prom_inst_1.INIT_RAM_1A = 256'h4105114411455FE180F55D9971FBE944B197EBCA253BAF0816F34EDA7E5A49CB;
defparam prom_inst_1.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF82A82882A88AA2A80001F5DD7400055405505;
defparam prom_inst_1.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_1.INIT_RAM_20 = 256'h89B6D9E53E438C2E51415405516FEFAB8040FFC13B5692820CDDDC2D141B6650;
defparam prom_inst_1.INIT_RAM_21 = 256'hA0013BE13E83F0C29C2718F4EAC5C9FE51015541412AFAFEB5107FC13ED3E0D7;
defparam prom_inst_1.INIT_RAM_22 = 256'h45051014405FBAAAF5156FE00BC2F1B6CC7778B5FBF488E155011550450BBBEF;
defparam prom_inst_1.INIT_RAM_23 = 256'hCA7673D7F17B671B45040005005BEEFEE4046EA40E90B1A3DF362192EAAC7385;
defparam prom_inst_1.INIT_RAM_24 = 256'hE4152AA05BC0F1F19327329F804A486E45540001114ABBEFB5113EB05ED5A1A4;
defparam prom_inst_1.INIT_RAM_25 = 256'h44501501450FAEFFB4006BB05B84E1A58366634F15079DB144500501410BAEAA;
defparam prom_inst_1.INIT_RAM_26 = 256'h26DB6794F90E30B84505501545BFBEAE0103FF04ED5A4A08337770B4506D9941;
defparam prom_inst_1.INIT_RAM_27 = 256'h8004EF84FA0FC30A709C63D3AB1727FA4405550504ABEBFAD441FF04FB4F835E;
defparam prom_inst_1.INIT_RAM_28 = 256'h14144051017EEAABD455BF802F0BC6DB31DDE2D7EFD2238454045541142EEFBE;
defparam prom_inst_1.INIT_RAM_29 = 256'h29D9CF5FC5ED9C6E14100014016FBBFB9011BA903A42C68F7CD8864BAAB1CE14;
defparam prom_inst_1.INIT_RAM_2A = 256'h9054AA816F03C7C64C9CCA7E012921BB15500004452AEFBED444FAC17B568693;
defparam prom_inst_1.INIT_RAM_2B = 256'h11405405143EBBFED001AEC16E1386960D998D3C541E76C411401405042EBAAB;
defparam prom_inst_1.INIT_RAM_2C = 256'h07E0ED6CE70D9E7D00004041411545501042BEBAED551AF85FB0A974E2388338;
defparam prom_inst_1.INIT_RAM_2D = 256'h4556ABEAE8504ABD13F52C29B78CDD3401405105505050055446ABFFBD555AAD;
defparam prom_inst_1.INIT_RAM_2E = 256'h15541450011544041116AABFA8410EE916F56939B79CD9650550111414410551;
defparam prom_inst_1.INIT_RAM_2F = 256'h07F5693965DD999315550441415011515016AAAAF8445EFC02E13828618989F3;
defparam prom_inst_1.INIT_RAM_30 = 256'h1542AFFEAC414AAD13F56828758DDD8255054445544544040446AEEBFC450EF8;
defparam prom_inst_1.INIT_RAM_31 = 256'h50005110011004015102AFBBF9501AB916E0394C65CD6DC65001410505145151;
defparam prom_inst_1.INIT_RAM_32 = 256'h1F83B5B39C3679F50001010504551540410AFAEBB5546BE17EC2A5D388E20CE1;
defparam prom_inst_1.INIT_RAM_33 = 256'h155AAFABA1412AF44FD4B0A6DE3374D30501441541414015511AAFFEF5556AB4;
defparam prom_inst_1.INIT_RAM_34 = 256'h5550514004551010445AAAFEA1043BA45BD5A4E6DE7365961540445051041545;
defparam prom_inst_1.INIT_RAM_35 = 256'h1FD5A4E59776664E5554110505404545405AAAABE1117BF00B84E0A1862627CF;
defparam prom_inst_1.INIT_RAM_36 = 256'h550ABFFAB1052AB44FD5A0A1D637760A5415111551151010111ABBAFF1143BE0;
defparam prom_inst_1.INIT_RAM_37 = 256'h4001444004401005440ABEEFE5406AE45B80E5319735B7184005041414514544;
defparam prom_inst_1.INIT_RAM_38 = 256'hFBEEBAEBBEFBEEBAC51451041145144104114510410451451041145144104114;
defparam prom_inst_1.INIT_RAM_39 = 256'h114510410451451041145144104514510EBAEFBEEBAEBBEFBEEBAEFBEFBAEBAE;
defparam prom_inst_1.INIT_RAM_3A = 256'h106FBEEBAEBBEFBEEBAEFBEFBAEBBEFBEEBAEBBEFBAEBAEFBE51041145144104;
defparam prom_inst_1.INIT_RAM_3B = 256'hBAEBBEFBAEBAEFBEFBA411451441045145104104514410411451441045145104;
defparam prom_inst_1.INIT_RAM_3C = 256'h104104514410411451441045145104114514EBAEBBEFBAEBAEFBEFBAEBBEFBEE;
defparam prom_inst_1.INIT_RAM_3D = 256'h14410EBBEFBAEBAEFBEFBAEBBEFBEEBAEFBEFBAEBAEFBEEBAEBBC51441045145;
defparam prom_inst_1.INIT_RAM_3E = 256'hBEFBAEBAEFBEEBAEBBEFBE410451451041145144104114510410451451041145;
defparam prom_inst_1.INIT_RAM_3F = 256'h145144104114510410451451041145144104516FBAEBAEFBEEBAEBBEFBEEBAEF;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[30:0],prom_inst_2_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 1;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'hFFFFFFFFFFD124A859628D444DA63848FDD7573FFFFFF48AA4F9FFFFFFFFFF03;
defparam prom_inst_2.INIT_RAM_01 = 256'h6073CE6F0F66538DDBBCCC96C1F27C20263200002100FB00126DB28053601615;
defparam prom_inst_2.INIT_RAM_02 = 256'hFFFFFFFFFFF9DA5E56A7D9BECCBDC0F2D64D425CCC82A0001DC42850216A4444;
defparam prom_inst_2.INIT_RAM_03 = 256'h7FBF963A6F77F37BBF3F77FDFAFDEBFBF6D85EFDAAAABFABAEFFD054545EBBAA;
defparam prom_inst_2.INIT_RAM_04 = 256'h2A76653E3282A9BDF075FBBFC0D172CA0FFDFF41D474187F374DFD4BF9BD4BF3;
defparam prom_inst_2.INIT_RAM_05 = 256'hF90BD43434343C20FA734343D4FEC6EF17788A72093926ED4BF5FB9F942FD3A3;
defparam prom_inst_2.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFF69BDCF77E8F9EFA894BDDF7BFDB17F7BFDFEE5FBF63F6E6E5;
defparam prom_inst_2.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC4B9E867A0973D096;
defparam prom_inst_2.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_0C = 256'h31131113322212A765976EDEDD26F6E9F169B78B3BDBAC19A3C488949DB6CA4B;
defparam prom_inst_2.INIT_RAM_0D = 256'h155BB14B6D8BA2A00E0072AB405DA016334486314CDB6AE66CB5732707531331;
defparam prom_inst_2.INIT_RAM_0E = 256'h5BCB2F345040CB540158556ED5D24B6E925B05050D558556EC011585A92B0056;
defparam prom_inst_2.INIT_RAM_0F = 256'h187E6C502A6A19F54640803484FD9085482627930013903EA4286D93EBAEB0F7;
defparam prom_inst_2.INIT_RAM_10 = 256'h8B800A40924BC452146D78F20AC489B4F404D9018C9630C5664116132D62524B;
defparam prom_inst_2.INIT_RAM_11 = 256'h0DF6CB3271DC60F9899B34D76C9CD21AB775935982278C948E07291A2AB6EF6A;
defparam prom_inst_2.INIT_RAM_12 = 256'hDFDEEA0FF9D5B1FB5364CEBFD7E40C8A2D5B565CCBDAD6BDFB5EE4937B5AFD55;
defparam prom_inst_2.INIT_RAM_13 = 256'hA836AD19BBAEABE06DC9949393252713224E26549C2449382452701324E00050;
defparam prom_inst_2.INIT_RAM_14 = 256'hBAC43C88D52CF466EEBAAC200046466EEBA5B466EEBA9610000000008F891231;
defparam prom_inst_2.INIT_RAM_15 = 256'hE028303D53AC96C9246D5F11BB95709564B6C51BE492CBCF75E5728DDC9B559B;
defparam prom_inst_2.INIT_RAM_16 = 256'hFFFFFFF5277E4D5555956C5B9359D936764D9326D922EBD92775F0DA601940E6;
defparam prom_inst_2.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_2.INIT_RAM_18 = 256'hD75DDDDD75FD5555F7DDD6A0A8A0AAA22A88175757F5EA082DD622205FF57DD4;
defparam prom_inst_2.INIT_RAM_19 = 256'h004E08A208A2208882222222222220888228820B7D7D7D7F55FFD55555FF57F5;
defparam prom_inst_2.INIT_RAM_1A = 256'h6402C93309983B040C947B2BD4CE0BC7ACB6122F9300530903066200004C6200;
defparam prom_inst_2.INIT_RAM_1B = 256'h000C0400040000926C02EC9433D0C804257614800D1349A4F64CA40D81480102;
defparam prom_inst_2.INIT_RAM_1C = 256'h24F1133292C8114E4B01B299C89120020005B6489644B8401209764B0200C000;
defparam prom_inst_2.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB8AC68A91236;
defparam prom_inst_2.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_2.INIT_RAM_20 = 256'hE855A1442B589750AAC4BA15589D42AC4E85589DB1D138D7CAC8000444554121;
defparam prom_inst_2.INIT_RAM_21 = 256'h21A8027883441C20D1070801B1029359AE324EA15685142B589D0AB50A215AC4;
defparam prom_inst_2.INIT_RAM_22 = 256'h6AC3804FF5600FF6ABFF5578F66BCF77E30790D0341B31E499F1B5DFDAAFC60F;
defparam prom_inst_2.INIT_RAM_23 = 256'hB5438277F14027F0B20A16917D70E0E1FE704EFE142D2F541EC01FE5270FE165;
defparam prom_inst_2.INIT_RAM_24 = 256'h914044EFE142D2EC8913B80003F9122780FECBC2C9C58C0180004FEC60080FE5;
defparam prom_inst_2.INIT_RAM_25 = 256'hDE3F79C78FDE394A5097B2280C0003BF9100409FC2C8285A5CBDB2200C01C03F;
defparam prom_inst_2.INIT_RAM_26 = 256'h1E50793D078F61E501E3D078E5294E4C94997C795E3B783D785E3B1E3979DE4F;
defparam prom_inst_2.INIT_RAM_27 = 256'hC88DABFF5CF8B267C931E30790D6823A5266D89E7078F41E0FC1E7078F4078FC;
defparam prom_inst_2.INIT_RAM_28 = 256'h949783B6D2F1DCF1DB264ADCF1DB29783978EDB6AFED35E3689F3D478C1E4358;
defparam prom_inst_2.INIT_RAM_29 = 256'h1DBE4C96F89E3B65A0F07B0F1DB29C2DE3B6D73C76F1E6CACBC71B6B78E5E4ED;
defparam prom_inst_2.INIT_RAM_2A = 256'hBE94A71D30F1DB2F89E3B878E36F83C79BA9878EC1E4ED95D8783B7DE0F1E80F;
defparam prom_inst_2.INIT_RAM_2B = 256'hDA5A5E0FDE3B77BC76EBC78EDDF3C76FA4D97D9E3B78E37DBC79BAB78EDF6F1D;
defparam prom_inst_2.INIT_RAM_2C = 256'h57DE39793B6CBC1DB2D78E36EBC79B294E52B78F478ED9A3C76DB5E0ED9AF276;
defparam prom_inst_2.INIT_RAM_2D = 256'h6F9878EDB4C4F1DB66278ED9793652E278FC1E38D9F0F1E6DBE1E3B67C3C76CA;
defparam prom_inst_2.INIT_RAM_2E = 256'h71BF41E3CDD4A4E52F878EC078EDD603C76FAC1E0EDD60F276FA52EC3C1C83C7;
defparam prom_inst_2.INIT_RAM_2F = 256'h05ECE48E23DC499742CE48E2FD71E52EB1C280BCF30F1EC3C1DBF41E4EDD6C3C;
defparam prom_inst_2.INIT_RAM_30 = 256'h2EB3263840902010160481205816DE0CF36E20CBA6F247869024080402204816;
defparam prom_inst_2.INIT_RAM_31 = 256'h65D00FE80100404020020080405A7393C832E80044A3C0CE4F24CBA0026571E5;
defparam prom_inst_2.INIT_RAM_32 = 256'h38835C5FA2B389E49AE2B47A0002008040400802010175E4F24CB8BD9C6F0712;
defparam prom_inst_2.INIT_RAM_33 = 256'h4816058101E3CE0E33CC29670719E6002017E90240B02C080440902C0B02F670;
defparam prom_inst_2.INIT_RAM_34 = 256'h1204022048160581204DCE4F3C932E81119C9E79265C22D28081205813020220;
defparam prom_inst_2.INIT_RAM_35 = 256'h10202010090E7071C41974C08E7279E49832E110240B02C0902026D204816058;
defparam prom_inst_2.INIT_RAM_36 = 256'h81008817F3838E20C997088ACE4F3C93065D02048160581207D6A02048160581;
defparam prom_inst_2.INIT_RAM_37 = 256'hE2CE4F3C93265C22F59C9E79260CBA6040902C0B024090202BD2048160581204;
defparam prom_inst_2.INIT_RAM_38 = 256'h832E911119C9E79260CBA6040902C0B02409025AD010240B02C0902204040201;
defparam prom_inst_2.INIT_RAM_39 = 256'hF220C99708881205816048120581015A90240B02C090240B02013026E7279E49;
defparam prom_inst_2.INIT_RAM_3A = 256'h816048120581F5280812058160481204C08080402C59C1C719264CB845E7393C;
defparam prom_inst_2.INIT_RAM_3B = 256'h0481605812048160581009815F3838E324C1974888BCE0E38C93065D35C81205;
defparam prom_inst_2.INIT_RAM_3C = 256'h20160CE4F3C8833265C22719C9E7910660CBA6040902C0B0240902C0B02022D2;
defparam prom_inst_2.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF90240B02C090240B02604040;
defparam prom_inst_2.INIT_RAM_3E = 256'h8E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38;
defparam prom_inst_2.INIT_RAM_3F = 256'hE38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E38E;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[30:0],prom_inst_3_dout[1]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 1;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h65B2C965B2472E72CADE68034004191B710D66805FEA87681100006200004021;
defparam prom_inst_3.INIT_RAM_01 = 256'hF0992F37511CC4473110CC4500C4DCCC4C44C42C4DCCC4C5478C04010165B2C9;
defparam prom_inst_3.INIT_RAM_02 = 256'h27BDA68EEA9764D347559B2EC4467E277ABB2EF6BDCA20113113313351100643;
defparam prom_inst_3.INIT_RAM_03 = 256'hCD0BEC8C881622672E31620E5F27326065F67326065F60A08165F20A0C165F27;
defparam prom_inst_3.INIT_RAM_04 = 256'h5060B2F937D8E7616FB61F67731D6062AA0C648A4C96D97639DB3CDD119BBBBE;
defparam prom_inst_3.INIT_RAM_05 = 256'h56DBD6473C00902D5CD54C55967922B220C0321400B3B35A3FAA732D966309F0;
defparam prom_inst_3.INIT_RAM_06 = 256'h0059FC0127D0049984DC00906E613705041B2FB17C9F320F305F4E4DC2ADB7A1;
defparam prom_inst_3.INIT_RAM_07 = 256'h95454800185EAEA7BDAD7DEC92200FCD67C79D7FD69A270094D338049F40127D;
defparam prom_inst_3.INIT_RAM_08 = 256'h3DCB879D9CB384FB7A23C76EECECEEA660296930AA669296930ACA2E4CA86A19;
defparam prom_inst_3.INIT_RAM_09 = 256'h94AFBE696D7BBA105400048024580AF63E002400039481018E35A726E7250802;
defparam prom_inst_3.INIT_RAM_0A = 256'hB5F5A972B657F25147A74016631EA2857D4702732C8B3641D2E2E8450EA9115F;
defparam prom_inst_3.INIT_RAM_0B = 256'hE4B01C705531333157570036FFB25B5240B2B6D929657F6E54A4B5F5B9720AEC;
defparam prom_inst_3.INIT_RAM_0C = 256'h1496848E5A19009251B196407020381141C0801009B04A0906E9B988C0508114;
defparam prom_inst_3.INIT_RAM_0D = 256'h6E692C6F474D352D6BE42D429A546B4D04928D8CB0238011C0980E0400804A59;
defparam prom_inst_3.INIT_RAM_0E = 256'hDF0E01E90C6BA798A5B2709011086C10EDB6C866DA5D232ED90CD96596596596;
defparam prom_inst_3.INIT_RAM_0F = 256'hBD50EE492492492408822AAC778F1E3EFBEFBF1F7E3F80FA262013635B7F1416;
defparam prom_inst_3.INIT_RAM_10 = 256'h96A00074A9522AA72BB44ED548B0096D5551A6CD48B0096D55402BB3000FF818;
defparam prom_inst_3.INIT_RAM_11 = 256'h19D77D242B1ED090C096ACDB8A7AB01B5A7CEDECE0CEBBA12158D68713500240;
defparam prom_inst_3.INIT_RAM_12 = 256'h16224D316BDA9B264C6CA6C9643A2F9557691B6EA3665585BB56037B4FFDBDFC;
defparam prom_inst_3.INIT_RAM_13 = 256'hD05BF82F82FC28C11214D9517C806B1DE8E89D42940014A457A3A5346BA2FC42;
defparam prom_inst_3.INIT_RAM_14 = 256'hAD51FCF924BE2B62705F8CA98CA796479257053C7DEE3B490AC17217242EC2E4;
defparam prom_inst_3.INIT_RAM_15 = 256'hB7492495FDB1B1E194A0F1B9E0F1BC4E3E87C078F87F4E3C9E5E3A7E17C36847;
defparam prom_inst_3.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF91DDCD080AED6F5FC3DF;
defparam prom_inst_3.INIT_RAM_17 = 256'h0000000000000000000000000000000000000BCF000103461E93000420155008;
defparam prom_inst_3.INIT_RAM_18 = 256'h0000FFFFFFFFFFFFFFFF000000000000FFFFFC00FFFFFFFFBA01FFFF00000000;
defparam prom_inst_3.INIT_RAM_19 = 256'h55555EBD55444155FEFFFFFFFEBFFA93FFFFFFFFFFEF5053FFFFFFFFEFAAAAAA;
defparam prom_inst_3.INIT_RAM_1A = 256'h405505410510E214017FFE716771C075F5609D03AF2D76AC3C9DB2DAF7740A76;
defparam prom_inst_3.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF8A208A02A82882A88AA2088001F5DD7400055;
defparam prom_inst_3.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_3.INIT_RAM_20 = 256'hD7A092CDF3D8F57E45100550404004416FAFBF9000FAD13B5392825C9DDC2C04;
defparam prom_inst_3.INIT_RAM_21 = 256'h4FEFEEE0017BA12B82A4C69C331CB4FE44501554510501401EBAFF80012EB13B;
defparam prom_inst_3.INIT_RAM_22 = 256'h54405015041514404EBAAAE0156FE44AC2A4F6CC726CF5BF4440555511155515;
defparam prom_inst_3.INIT_RAM_23 = 256'hD0E4A5CB3337D6E154414005445005410BFEFEE4142AF45E90F0A3DF762093BA;
defparam prom_inst_3.INIT_RAM_24 = 256'h1BEEAFB4116AE05AC0B5B1937337DB8014410001404541154EBFEFF4153BB45E;
defparam prom_inst_3.INIT_RAM_25 = 256'h11440054511505454EAEFAA4113BA04B80A1A4C722660F111145004151155040;
defparam prom_inst_3.INIT_RAM_26 = 256'h5E824B37CF63D5F81440154101001105BEBEFE4003EB44ED4E4A09727770B010;
defparam prom_inst_3.INIT_RAM_27 = 256'h3FBFBB8005EE84AE0A931A70CC72D3FA11405551441405007AEBFE0004BAC4EF;
defparam prom_inst_3.INIT_RAM_28 = 256'h51014054105451013AEAAB8055BF912B0A93DB31C9B3D6FF1101555444555455;
defparam prom_inst_3.INIT_RAM_29 = 256'h4392972CCCDF5B8551050015114015042FFBFB9050ABD17A43C28F7DD8824EEA;
defparam prom_inst_3.INIT_RAM_2A = 256'h6FBABED045AB816B02D6C64DCCDF6E0151040005011504553AFFBFD054EED17B;
defparam prom_inst_3.INIT_RAM_2B = 256'h45100151445415153ABBEA9044EE812E0286931C89983C444514010544554100;
defparam prom_inst_3.INIT_RAM_2C = 256'h501AA807E1ED78A311110501405105511545500003EBBAED550AF80BF0B975E2;
defparam prom_inst_3.INIT_RAM_2D = 256'h0545514556EBAAFD415BBD13F12828A710511405501115544010041043EBEFBD;
defparam prom_inst_3.INIT_RAM_2E = 256'h04451055550450011450040516EABFE9450BE907E56939F21441141554101005;
defparam prom_inst_3.INIT_RAM_2F = 256'h411FB816B17C396404441054154441504005515016EEEAA8445FFC02A1392870;
defparam prom_inst_3.INIT_RAM_30 = 256'h1011540546EFBEAC504FAD13A56D287544445050014105544540004416EFEFFC;
defparam prom_inst_3.INIT_RAM_31 = 256'h44444140005110004104015142FFABE8541AB916A13C09614444515000511405;
defparam prom_inst_3.INIT_RAM_32 = 256'h406AA01F87B5E28D4444140501441544551540000FAEEBB5542BE02FC2E5D789;
defparam prom_inst_3.INIT_RAM_33 = 256'h151545155BAEABF5056EF44FC4A0A29F4144501540445551004010410FAFBEF5;
defparam prom_inst_3.INIT_RAM_34 = 256'h1114415554114004514010145BAAFFA5142FA41F95A4E7CA5104505550404014;
defparam prom_inst_3.INIT_RAM_35 = 256'h047EE05AC5F0E5931110415055110541001545405BBBAAA1117FF00A84E4A1C2;
defparam prom_inst_3.INIT_RAM_36 = 256'h404550151BBEFAB1413EB44E95B4A1D61111414005041551150001105BBFBFF1;
defparam prom_inst_3.INIT_RAM_37 = 256'h1111050001444001041005450BFEAFA1506AE45A84F025871111454001445014;
defparam prom_inst_3.INIT_RAM_38 = 256'h4514514504104104145145145041041041051451451410410410514514514504;
defparam prom_inst_3.INIT_RAM_39 = 256'hFAEBAEBAEBEFBEFBEFAEBAEBAEBEFBEFB4514104104105145145141041041041;
defparam prom_inst_3.INIT_RAM_3A = 256'h043EFBEFBEFAEBAEBAEBEFBEFBEFAEBAEBAEBAFBEFBEFBEBAEBAEBAFBEFBEFBE;
defparam prom_inst_3.INIT_RAM_3B = 256'h5145041041041451451450410410414514514514104104105145145141041041;
defparam prom_inst_3.INIT_RAM_3C = 256'hAEBAEBEFBEFBEFAEBAEBAEBEFBEFBEFAEBAE1041051451451410410410514514;
defparam prom_inst_3.INIT_RAM_3D = 256'h51451EFAEBAEBAEBEFBEFBEFAEBAEBAEBEFBEFBEFBEBAEBAEBAFBEFBEFBEBAEB;
defparam prom_inst_3.INIT_RAM_3E = 256'h0410410414514514504104104145145145041041041051451451410410410514;
defparam prom_inst_3.INIT_RAM_3F = 256'hFBEFBEFBEFAEBAEBAEBEFBEFBEFAEBAEBAEBEF94514514104104105145145141;

pROM prom_inst_4 (
    .DO({prom_inst_4_dout_w[30:0],prom_inst_4_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_4.READ_MODE = 1'b0;
defparam prom_inst_4.BIT_WIDTH = 1;
defparam prom_inst_4.RESET_MODE = "SYNC";
defparam prom_inst_4.INIT_RAM_00 = 256'hFFFFFFFFFFD861867D004E594C6CF201FD1898BFFFFF80555EF8FFFFFFFFFF90;
defparam prom_inst_4.INIT_RAM_01 = 256'h206BCC680621438D9F300404C1D0352015260000E002CC000A63748142C33C4F;
defparam prom_inst_4.INIT_RAM_02 = 256'hFFFFFFFFFFFA0CA06783E9F68C895EB35551A58B00496FF002276EDDB951FFFF;
defparam prom_inst_4.INIT_RAM_03 = 256'h77C2A97A6AD85356C27AD85E1056415CBFF8650A0020AB830AAAFFFAFFF00105;
defparam prom_inst_4.INIT_RAM_04 = 256'h35B046D923034EC8802616CA0120A9E68FAE16A7ADEB7885774D7A9C29AA9C27;
defparam prom_inst_4.INIT_RAM_05 = 256'h16F40A4A4A4A4BDD02A226258DC5BD10288142A29A5A570A9C2214312B70AC82;
defparam prom_inst_4.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFC0CA35A58F2D4BCF084A028B155B849412156E146A6254D4E;
defparam prom_inst_4.INIT_RAM_07 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_4.INIT_RAM_08 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_4.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD00D7EF7FA01BFC00;
defparam prom_inst_4.INIT_RAM_0A = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_4.INIT_RAM_0B = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_4.INIT_RAM_0C = 256'h9999BB9BB9E24003000A906DC4836E2422966114CDB89066608A4C0049DA0200;
defparam prom_inst_4.INIT_RAM_0D = 256'h2810DF07F6F8F3DB36B285217086C3151340B42D8D8C8E46CE4767738DD99B99;
defparam prom_inst_4.INIT_RAM_0E = 256'hD8A34335B148EFD9FE28A047F73FFDB9FFEDDF5F47A28A047E7E62811FD0D98A;
defparam prom_inst_4.INIT_RAM_0F = 256'hC752A0A96AAF1AB7C6BD2AB50074DDF49D226581B00106A800014C01966E8ACC;
defparam prom_inst_4.INIT_RAM_10 = 256'hC2DB6DB2DD3ECA69956B4860E4A9208068DF6D11C7BBF20D42408E4141453443;
defparam prom_inst_4.INIT_RAM_11 = 256'h9464801010C4696AA0080555680C5116A55542C42383460F8783F6EC45DB6FF3;
defparam prom_inst_4.INIT_RAM_12 = 256'hD7DEE0ED7DDF81F849B689C05FF6E669761D87FEFC6718C61CE71B6D8CEBFF5C;
defparam prom_inst_4.INIT_RAM_13 = 256'h7627E80CEECBFA308A20AB78415AF0815DE102ABC200B78400AF08005E100014;
defparam prom_inst_4.INIT_RAM_14 = 256'hEC901E8EFFA96033BB2FE8115518033BB2F56033BB2FD408AAAAAAAA36909219;
defparam prom_inst_4.INIT_RAM_15 = 256'hC86433F4FE9FFBFDBF973B9045FB3A05FEBB6BA8F52D34349A988D48C8C860CE;
defparam prom_inst_4.INIT_RAM_16 = 256'hFFFFFF84827F54AAAA2A80A82869AAD66AB7ADDAD936F34ADED32EEEF4FDFDDF;
defparam prom_inst_4.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_4.INIT_RAM_18 = 256'hA28A0A0A80AAAAAAA02821DDDF7F555F5DF555DD55D560888AA000002228A880;
defparam prom_inst_4.INIT_RAM_19 = 256'h0A6A02A0A80A0A8280A0A0A0A0A0A2828A08208208A208A22288888888882228;
defparam prom_inst_4.INIT_RAM_1A = 256'h00628408C01DBA62800C40351EEA5043A284101001B001806A8200800A680080;
defparam prom_inst_4.INIT_RAM_1B = 256'h1C4AE5EAA1C1EFFADAD9FED96890447510FFB1C0FB8EE336BF0408FFD542AC05;
defparam prom_inst_4.INIT_RAM_1C = 256'h007080018D06788207C811CD6EDDF150F3F7FB6DFB51455C5BE2FF02A0E2BCAA;
defparam prom_inst_4.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF94022476DBCB;
defparam prom_inst_4.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_4.INIT_RAM_20 = 256'h729DCA694B592BA54AC95CA9592E94AC9729592EBAD258F6C356000110004570;
defparam prom_inst_4.INIT_RAM_21 = 256'hF804E04F127895C4AE24F10E6E209059EE24974A7729A94B592E53BA534A5AC9;
defparam prom_inst_4.INIT_RAM_22 = 256'h90542A96A82AB6B367293B106DD8B6EE411D7C0AEDF4EC53772042210114823A;
defparam prom_inst_4.INIT_RAM_23 = 256'h40142A9B58154B563362C69842050136D405536AC58D3480A5556D6029B6AD26;
defparam prom_inst_4.INIT_RAM_24 = 256'hC45D5936AC58D3532164EAEAEDAE42C9BB6B029A4F5B25760E8E96B923A3B6A1;
defparam prom_inst_4.INIT_RAM_25 = 256'h265C9929972659084B056CC3B87474DAE61D1D2D58CD8B1A682B6883B0B24EDA;
defparam prom_inst_4.INIT_RAM_26 = 256'hE663995C39978E64B265EB996421280090019299265C985C99265C265C992657;
defparam prom_inst_4.INIT_RAM_27 = 256'hBCE94420A21001108088411D7C02E0FC40074B264B9970E6572E663997AC9978;
defparam prom_inst_4.INIT_RAM_28 = 256'h852995D69532D132E900429132EB0A985A9974C99CA6EE409762CA310475F00B;
defparam prom_inst_4.INIT_RAM_29 = 256'h2E94008523A65D691730B5732E90864265D6954CB532CA4294CB2B48996A6574;
defparam prom_inst_4.INIT_RAM_2A = 256'hB08421925732EB4AB2658B9975215CCB2B4AB9960E65748403985D695732D593;
defparam prom_inst_4.INIT_RAM_2B = 256'hF215A656A65D214CBAD2A9974854CBAC200850265E9965234CB2B4C9974A932E;
defparam prom_inst_4.INIT_RAM_2C = 256'h18A65E985D334CAEBC89975384CBAB884218699629974C14CBAE2A6174E530BA;
defparam prom_inst_4.INIT_RAM_2D = 256'hA64B9975C61D32E992C9975C7002190E9978E6594ED732EAE30E65D325CCBAE2;
defparam prom_inst_4.INIT_RAM_2E = 256'hB29D2E65D5E43021A639970E9974C964CBAF38E6574ED730BAE219B5CCAE5CCB;
defparam prom_inst_4.INIT_RAM_2F = 256'h93336156452CBAFF9A365176D0475F0A2D70083A49732F1CC2E99AE6575C65CC;
defparam prom_inst_4.INIT_RAM_30 = 256'h020EF18E721C8E464390E4390E4426117257597FE5328B241C872392C9390E43;
defparam prom_inst_4.INIT_RAM_31 = 256'hBFF32203E479192C97C8F23919144D85D75FF3392145D03617597FCCC948075F;
defparam prom_inst_4.INIT_RAM_32 = 256'h5D657C80560DE2EB2BF6410027C8F239191F23C8E464026565D7FE02AE132B2E;
defparam prom_inst_4.INIT_RAM_33 = 256'h0E4390E4641136175595109B0BAAC8CC964A41C8721C872592721C8721C909BC;
defparam prom_inst_4.INIT_RAM_34 = 256'h4792C9390E4390E4793A36175975FF36266CACBACBFF698C08E4390E49C8C939;
defparam prom_inst_4.INIT_RAM_35 = 256'hBC8C964B26D1B2B2EB2FF95219B0BACBAF5FF21C8721C8723C8C990390E4390E;
defparam prom_inst_4.INIT_RAM_36 = 256'hE4B25E4E8D9597597AFF931336175975EBFE6390E4390E47936302390E4390E4;
defparam prom_inst_4.INIT_RAM_37 = 256'hDA36565D65EBFE56D46CACBACB97FCA8721C8721C8F23C8C998390E4390E4791;
defparam prom_inst_4.INIT_RAM_38 = 256'hE5FF2B6B26CACBACB97FC8C721C8721C8F23C890811C8721C8723C979192C964;
defparam prom_inst_4.INIT_RAM_39 = 256'h65597AFF958E4390E4391E4791E464841C8721C8723C8F23C964BC949B2B2EB2;
defparam prom_inst_4.INIT_RAM_3A = 256'hE4391E4791E400C08E4390E4391E4792F232592C8306C2EB22EB97FE8884D85D;
defparam prom_inst_4.INIT_RAM_3B = 256'h90E4390E4791E4791E4B25E484D85D645D7AFFD1311361759175EBFF428E4390;
defparam prom_inst_4.INIT_RAM_3C = 256'h9649B3617595645EBFE56966CACBA2EABD7FE8C721C8721C8F23C8F23C8C9D03;
defparam prom_inst_4.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9C8721C8723C8F23C979192C;
defparam prom_inst_4.INIT_RAM_3E = 256'h0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0;
defparam prom_inst_4.INIT_RAM_3F = 256'hFC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0FC0F;

pROM prom_inst_5 (
    .DO({prom_inst_5_dout_w[30:0],prom_inst_5_dout[2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_5.READ_MODE = 1'b0;
defparam prom_inst_5.BIT_WIDTH = 1;
defparam prom_inst_5.RESET_MODE = "SYNC";
defparam prom_inst_5.INIT_RAM_00 = 256'h0100904824860A149216E8074024120DA501EE800AFF850D097FFFE2FFFF400E;
defparam prom_inst_5.INIT_RAM_01 = 256'h00D2413BB9AEEE6BFF9AEEE73266FEE66E66CC866FEE66E733CDA602C8482402;
defparam prom_inst_5.INIT_RAM_02 = 256'h0830196319A1020CB8CD2810066083304202300AC00C283B99B999BBF99B61B8;
defparam prom_inst_5.INIT_RAM_03 = 256'h69AC08440000191270100083600520483604520483604190CA4604190CA46048;
defparam prom_inst_5.INIT_RAM_04 = 256'hC865230228114B4150242048522CF933990CBD522004801018522EA160EAA4A8;
defparam prom_inst_5.INIT_RAM_05 = 256'h7B6DD46804DBFCFFF6776EF6FB0FB0DB176D80937C044CC3412E420800221230;
defparam prom_inst_5.INIT_RAM_06 = 256'hBE0E06F8783BE1517460DBFCDC5D180C865230208023216BAE2302010EF6DBA7;
defparam prom_inst_5.INIT_RAM_07 = 256'hC864B65B67EBCF918D634EA6FB812D454E9D3E26132CB87C19E7C3E0E06F8381;
defparam prom_inst_5.INIT_RAM_08 = 256'h1E12F5A1201C238A8E328862E101033776E5E1A6F3776E5E1A6F7DF368F0899D;
defparam prom_inst_5.INIT_RAM_09 = 256'h84DA8C49247B3F044926DB650AD89C4146139B2DB04C31FD24988100810CC090;
defparam prom_inst_5.INIT_RAM_0A = 256'h7A4EFDDB49E91B68E00804F4BBA00FD680079E503C4F006173E0E98FAB271352;
defparam prom_inst_5.INIT_RAM_0B = 256'h207C44B5CCB9BB99FFDD96C9005B7FAFD3497FFFF69E91BB76D25A46FDFBADBB;
defparam prom_inst_5.INIT_RAM_0C = 256'hC28B0331ED86627BB44AAC20021001D628008D150F2569A50002062B11906788;
defparam prom_inst_5.INIT_RAM_0D = 256'h26BD539038D888017C9BD23DB1200BF613DDA355432011900EB3400468A87184;
defparam prom_inst_5.INIT_RAM_0E = 256'hFD8C1C4A12AAA22869803C023C98A39965064CA2825505AA50848C30C30C30C3;
defparam prom_inst_5.INIT_RAM_0F = 256'hDDF074000000000001405552004081000000008001018EDB02737DB3FFFF103F;
defparam prom_inst_5.INIT_RAM_10 = 256'h4F986DD89F2D864786D8CFE52DD9BE9320C3836D2DD9BE9320C206DB36CDFC8F;
defparam prom_inst_5.INIT_RAM_11 = 256'h8CE326F73FDB9D6C30DEBA6DE963791B7E79487974671937B9FEDCE7B9CB6DB3;
defparam prom_inst_5.INIT_RAM_12 = 256'h14134111FFDA4DB44222936FB4C23F9DD7F10DEB99B45AD7246F226FCF090F0E;
defparam prom_inst_5.INIT_RAM_13 = 256'h4D734EBAEBB724AD1A126DD0BCDA29F766A5C0E08EE7F5E7DD9A94B20A043672;
defparam prom_inst_5.INIT_RAM_14 = 256'h21810081120081627C5A5BA75A999469D85E084F9FF3CFCE4BF5D55D5ABAABAB;
defparam prom_inst_5.INIT_RAM_15 = 256'h4D8B6C90AF2323621A6DFBABE2E1B84E39AF2578E49C92180C1624F9B6C3F884;
defparam prom_inst_5.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA426D80109356C0AC420;
defparam prom_inst_5.INIT_RAM_17 = 256'h00000000000000000000FFFFFFFFFFFF00000FD0000002C07E4D540905CBA740;
defparam prom_inst_5.INIT_RAM_18 = 256'h0000000000000000000000000000000000000020000103E7FBFE000000000000;
defparam prom_inst_5.INIT_RAM_19 = 256'hFFFFFEEFAAAFEBEFA4A2AAAA94420500AAAAAAAABA9A0502AAAAAAAA713FFFFF;
defparam prom_inst_5.INIT_RAM_1A = 256'h400055405500A210C2DB33854061803457E49529037D56248A96DA48F67F1358;
defparam prom_inst_5.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFAA08288A208A02A82882A80AA2088001F5DD7;
defparam prom_inst_5.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_5.INIT_RAM_20 = 256'h2BB17BD7A597D9A604140405510015005044417FAAEF9050AEC13A0792925C8D;
defparam prom_inst_5.INIT_RAM_21 = 256'h5005144FAFBEE0006BE02B83A5C2C92304541541400504545505416FAFEAF005;
defparam prom_inst_5.INIT_RAM_22 = 256'h10505554404051000500404FBAEBE0557BB04BD3B1E6DD770054555044145140;
defparam prom_inst_5.INIT_RAM_23 = 256'h3AA41EC1E4F0DA2210515555000014551011410BBEFEA0402AF44E90B1A3DF27;
defparam prom_inst_5.INIT_RAM_24 = 256'h1010454FEEEEF4147BB51AC0E0B4867310015555110545404505110FEFAAF045;
defparam prom_inst_5.INIT_RAM_25 = 256'h11054001441054504505405FEEEAA4102BE05A80A4E0C2621105501540145100;
defparam prom_inst_5.INIT_RAM_26 = 256'hAEC5EF5E965F669B1050101544005401411105FEABBE4142BB04E81E4A497236;
defparam prom_inst_5.INIT_RAM_27 = 256'h4014513EBEFB8001AF80AE0E970B248C1150550500141151541505BEBFABC014;
defparam prom_inst_5.INIT_RAM_28 = 256'h41415551010144001401013EEBAF8155EEC12F4EC79B75DD0151554110514501;
defparam prom_inst_5.INIT_RAM_29 = 256'hEA907B0793C3688841455554000051544045042EFBFA8100ABD13A42C68F7C9D;
defparam prom_inst_5.INIT_RAM_2A = 256'h4041153FBBBBD051EED46B0382D219CC40055554441515011414443FBEABC114;
defparam prom_inst_5.INIT_RAM_2B = 256'h44150005104151411415017FBBAA9040AF816A02938309894415405500514400;
defparam prom_inst_5.INIT_RAM_2C = 256'hEBEFBD501BA817E150504110511405505105511544110003EBBAED554AE80AF0;
defparam prom_inst_5.INIT_RAM_2D = 256'h1450050545114543EABBFD415BBD13F150105114411415541115544011441043;
defparam prom_inst_5.INIT_RAM_2E = 256'h54145144441055550440011050440557EEBEE9440BE907A55410510445141555;
defparam prom_inst_5.INIT_RAM_2F = 256'hEFFEFC511FAC16B154145144445054054445504005151016EEEBA8445FFD02B1;
defparam prom_inst_5.INIT_RAM_30 = 256'h5114011015140546FFBBAC504FA813A514141144445150014105540550414016;
defparam prom_inst_5.INIT_RAM_31 = 256'h14141044444140001010004144515142FBABE8541BBD17A11414104444414000;
defparam prom_inst_5.INIT_RAM_32 = 256'hAFBEF5406EA05F864141044144501541441544551044000FAEEBB5552BA02BC3;
defparam prom_inst_5.INIT_RAM_33 = 256'h514014151445150FAAEFF5056EF44FC54041445104505550445551004510410F;
defparam prom_inst_5.INIT_RAM_34 = 256'h5051451110415554110004414110155FBAFBA5102FA41E955041441114505554;
defparam prom_inst_5.INIT_RAM_35 = 256'hBFFBF1447EB05AC55051451111415015111541001454405BBBAEA1117FF40AC4;
defparam prom_inst_5.INIT_RAM_36 = 256'h445004405450151BFEEEB1413EA04E955050451111454005041550154105005B;
defparam prom_inst_5.INIT_RAM_37 = 256'h5050411111050000404001051145450BEEAFA1506EF45E845050411111050001;
defparam prom_inst_5.INIT_RAM_38 = 256'h5145145145145145104104104104104104114514514514514514410410410410;
defparam prom_inst_5.INIT_RAM_39 = 256'h1451451451041041041041041045145145145145145144104104104104104104;
defparam prom_inst_5.INIT_RAM_3A = 256'hEF90410410410410410451451451451451451441041041041041041145145145;
defparam prom_inst_5.INIT_RAM_3B = 256'hEBAEBAEBAEBAEFBEFBEFBEFBEFBEFBAEBAEBAEBAEBAEBAEBBEFBEFBEFBEFBEFB;
defparam prom_inst_5.INIT_RAM_3C = 256'hBAEBAEFBEFBEFBEFBEFBEFBAEBAEBAEBAEBAEBAEBBEFBEFBEFBEFBEFBEEBAEBA;
defparam prom_inst_5.INIT_RAM_3D = 256'h14514FBEFBEFBEFBAEBAEBAEBAEBAEBAEFBEFBEFBEFBEFBEFBEEBAEBAEBAEBAE;
defparam prom_inst_5.INIT_RAM_3E = 256'h4514514510410410410410410451451451451451451441041041041041041145;
defparam prom_inst_5.INIT_RAM_3F = 256'h4104104104104104104514514514514514510410410410410410411451451451;

pROM prom_inst_6 (
    .DO({prom_inst_6_dout_w[30:0],prom_inst_6_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_6.READ_MODE = 1'b0;
defparam prom_inst_6.BIT_WIDTH = 1;
defparam prom_inst_6.RESET_MODE = "SYNC";
defparam prom_inst_6.INIT_RAM_00 = 256'hFFFFFFFFFFD041F2C00430404E0C1326FC64E4BFFFFFAEBAADF8FFFFFFFFFF44;
defparam prom_inst_6.INIT_RAM_01 = 256'hE392E24A83E5430D9FF4660EC3E335201356AAAAA050480002701860AAC69444;
defparam prom_inst_6.INIT_RAM_02 = 256'hFFFFFFFFFFFEA3871C824B706AA85C36C28B410B053C400508A7CFDF3C41BBBB;
defparam prom_inst_6.INIT_RAM_03 = 256'hC00AE960426152130A6261505504541880004428001011410045101044401504;
defparam prom_inst_6.INIT_RAM_04 = 256'h88B6715B38D08339202C52B8802930808038549525485015EC080258A90210AE;
defparam prom_inst_6.INIT_RAM_05 = 256'h52D4612321232F5409B48694A5D4B503981CC9B51D4C563218A05075696285B3;
defparam prom_inst_6.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFF008834A14624430600080A09504B141050510C50486A10D28;
defparam prom_inst_6.INIT_RAM_07 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_6.INIT_RAM_08 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_6.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF015F395CE02AE603;
defparam prom_inst_6.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_0C = 256'hAA88888AAA804383492F7146B5DA35AE79AA5BCCE8D6B86245E72E9074E4D901;
defparam prom_inst_6.INIT_RAM_0D = 256'hF74F7984BBCEF9C92C22A58030973DD59212112DBAFB8D77DDC6BBEFDCCAA8AA;
defparam prom_inst_6.INIT_RAM_0E = 256'h89216E9197583CB9275FDD397B0F3CF95D75BE7F3F35FDD3965B75F4F7EF6DD7;
defparam prom_inst_6.INIT_RAM_0F = 256'h4B5846B940CE91272449AA91A066CC4DE7046799A0414AB6069565C1AA471A66;
defparam prom_inst_6.INIT_RAM_10 = 256'hC7C9BC9BD9A5A14DD36D6CF0976D20A0524D2E31C52F029A6AD2B0410670A209;
defparam prom_inst_6.INIT_RAM_11 = 256'hD0C48010105569CB480A34A62008E25535499055E28346170B859273FA4BE8B1;
defparam prom_inst_6.INIT_RAM_12 = 256'hF2DE429D289C3C939EFAAC60161F223BB62D8B6AB6B5AD6B06318924C632C2BD;
defparam prom_inst_6.INIT_RAM_13 = 256'hDD530F2ECCEB13DC0E9D74B53AE56A7AE2D4F5D5A977CB5277D6A43BED4800FF;
defparam prom_inst_6.INIT_RAM_14 = 256'hCED00BAD3BEC6CBB33AC4C195500CBB33AC1BCBB33AC4604AAAAAAAA027846BA;
defparam prom_inst_6.INIT_RAM_15 = 256'h0ACC4249C8B3CF3EF37F6BEDE65C5E09D669609911C4105144A8146FBFAB5EEC;
defparam prom_inst_6.INIT_RAM_16 = 256'hFFFFFFA982711AAAAA6AB5A7E56A2AD28AB5AD5ACA76DBAA4816D236D4BDEA7F;
defparam prom_inst_6.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_6.INIT_RAM_18 = 256'h20822882228888888220820A0A800000A822220AAA88957F575C00002282A2A8;
defparam prom_inst_6.INIT_RAM_19 = 256'h0410000AA800AA802AA00AA00AA00A802A02A02A02A0A80A0A82828282820A08;
defparam prom_inst_6.INIT_RAM_1A = 256'h03BACC2D4058B3A7C0681D8972A840498C3E030219A04114AB1C390004103900;
defparam prom_inst_6.INIT_RAM_1B = 256'h5D66E1AAA1E5F0C8924D32CC67D2147150994B719A9FA3961908A9F6450AA801;
defparam prom_inst_6.INIT_RAM_1C = 256'h005888939DB99EF27514092566C9F1564BDE592E4B1CE35C59E29909A6EA68AA;
defparam prom_inst_6.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC6AE2C126FFF;
defparam prom_inst_6.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_6.INIT_RAM_20 = 256'h57B35EDBD9746AAF5BA355EB746ABDBA357B746A72A8D7B207C9000404454005;
defparam prom_inst_6.INIT_RAM_21 = 256'hF777FB5F2AB953CA9E54F2D3FE545ABF6570355ECD7B6BD9746AF66AF6DECBA3;
defparam prom_inst_6.INIT_RAM_22 = 256'h89142EF4C48BB4C8CD906ECAA37651B92A6FFBA77FD19920DD9106ECA33644DF;
defparam prom_inst_6.INIT_RAM_23 = 256'h44152D9A64177A6FA7FBF43F53054F369905F34DF7E87041E41769B079B4DDCE;
defparam prom_inst_6.INIT_RAM_24 = 256'h107DBF34DF7E876083ECA1EDED3107D97B4CBAFB9D6181F41EDEF4CC0FB7B4DD;
defparam prom_inst_6.INIT_RAM_25 = 256'h64D092D934E4D5EF7075A607A0F6ECD3303DBDE9BE9FEFD0EFAD2207A17E5ED3;
defparam prom_inst_6.INIT_RAM_26 = 256'hE4BF93D3F934BE4BF64D1F9357BDC1F8DFF1499264D192D092E4D3E4D29264F4;
defparam prom_inst_6.INIT_RAM_27 = 256'hFD7BEE997748CBBE67DD226FFBB97B257FC527E4979347E4F43E4BF934FD9349;
defparam prom_inst_6.INIT_RAM_28 = 256'hF7593D4FED26B326A7FC7BBF26A7F493D49353EFBE75DF2B3FE99774A9BFEEE5;
defparam prom_inst_6.INIT_RAM_29 = 256'h6A79F8F77FE4D4F68F25ADF26A7EF49E4D4F6DC9AD2699FBBC9A67B6935A4F53;
defparam prom_inst_6.INIT_RAM_2A = 256'h7B77BD26EF26A7B67E4D67934CFBBC9A67B67935BE4F53F75F92D4F6CF26B7B2;
defparam prom_inst_6.INIT_RAM_2B = 256'hEDDDA4F564D4F2C9A9FD59353CBC9A9FDF8F64E4D5934CFAC9AE7B59353CB26A;
defparam prom_inst_6.INIT_RAM_2C = 256'hD924D793D4FBC96A7B7934CF3C9AE7B77BD7493559353CBC9A9FDE4B53EF27A9;
defparam prom_inst_6.INIT_RAM_2D = 256'h9E779353FAFF26A7D5F9353DB7E3D9BF935FE4D73CEF2699FD7E4D4FABC9A9ED;
defparam prom_inst_6.INIT_RAM_2E = 256'hA67D7E4D73DBB3BD667935FF9353EEFC9A9FDDE4F53EFF27A9EDD9B3C96BFC9A;
defparam prom_inst_6.INIT_RAM_2F = 256'hFF336F34D1ABB6ADFE36F74DDD6BFFED35B2A3BA4CF26BFC9EA7DDE4B53DAFC9;
defparam prom_inst_6.INIT_RAM_30 = 256'hE517F2973FCFF7FFF9FE7F9FE7F0A6B74815DF56F1359AF2CFF3FDFFFF9FE7F9;
defparam prom_inst_6.INIT_RAM_31 = 256'hAB6FFA0C7F9FFFFFF8FF3FDFFFC72DAD76D5BFDFE85D74B6B5DF56DBFF412BFF;
defparam prom_inst_6.INIT_RAM_32 = 256'hD77D73E15F0DB6BBEB9F455A88FF3FDFFFE3FCFF7FFF0E6F5DB56F0269337AED;
defparam prom_inst_6.INIT_RAM_33 = 256'hE7F9FE7FFF5DB6F4DD73C25B5AE69BFFFFFA0CFF3FCFF3FFFF3FCFF3FCFF01B6;
defparam prom_inst_6.INIT_RAM_34 = 256'hF9FFFF9FE7F9FE7F9FE836B5D76D5BFEFA6DEBA6DAB6D052A27F9FE7FCFFFF9F;
defparam prom_inst_6.INIT_RAM_35 = 256'hCFFFFFFFFAE5B5A6BBEADF3D25B7A69BEBD5B6CFF3FCFF3FCFFFF099FE7F9FE7;
defparam prom_inst_6.INIT_RAM_36 = 256'h7FFFE7FA4DAD35DF56ADFF7D36F4D37D7AB6D9FE7F9FE7F9FC14A89FE7F9FE7F;
defparam prom_inst_6.INIT_RAM_37 = 256'h1CB6F5D36D7AB6DF096D69AEFAF56F9F3FCFF3FCFF3FCFFFF099FE7F9FE7F9FE;
defparam prom_inst_6.INIT_RAM_38 = 256'hAD5B6FEFC6D69AEFAF56FBF3FCFF3FCFF3FCFF2BD44FF3FCFF3FCFF9FFFFFFFF;
defparam prom_inst_6.INIT_RAM_39 = 256'h5CDB5EADB7E7F9FE7F9FE7F9FE7FFFECCFF3FCFF3FCFF3FCFFFFCFF91B7AE9B6;
defparam prom_inst_6.INIT_RAM_3A = 256'h7F9FE7F9FE7FD5AA27F9FE7F9FE7F9FF3FFFFFFFFBF6DE9A6EDAB56D9BBADAD7;
defparam prom_inst_6.INIT_RAM_3B = 256'hFE7F9FE7F9FE7F9FE7FFFE7FECDBD34DDB56ADB373636B5D737D7AB7D7E7F9FE;
defparam prom_inst_6.INIT_RAM_3C = 256'hFFFDFB6B5D736DD5AB7CD9D6DEBA66F9AB56D9B3FCFF3FCFF3FCFF3FCFFFFD19;
defparam prom_inst_6.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFF3FCFF3FCFF3FCFF9FFFFF;
defparam prom_inst_6.INIT_RAM_3E = 256'hF000FFF000FFF000FFF000FFF000FFF000FFF000FFF000FFF000FFF000FFF000;
defparam prom_inst_6.INIT_RAM_3F = 256'hFFF000FFF000FFF000FFF000FFF000FFF000FFF000FFF000FFF000FFF000FFF0;

pROM prom_inst_7 (
    .DO({prom_inst_7_dout_w[30:0],prom_inst_7_dout[3]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_7.READ_MODE = 1'b0;
defparam prom_inst_7.BIT_WIDTH = 1;
defparam prom_inst_7.RESET_MODE = "SYNC";
defparam prom_inst_7.INIT_RAM_00 = 256'h4100020925C32A100216C126402412049400AC00A0EA854F810000420000003E;
defparam prom_inst_7.INIT_RAM_01 = 256'h9052010888E33238888E222226AABA222A230DAAABA222A36859222288400092;
defparam prom_inst_7.INIT_RAM_02 = 256'h309659621D136F2CB0E9B934155312BB52D78A4A2AE3188888AAAAAAC8A9249A;
defparam prom_inst_7.INIT_RAM_03 = 256'hE1E88040D0A35D38635A35E58471831E58431831E5843B31085443B310854430;
defparam prom_inst_7.INIT_RAM_04 = 256'h98842A21810C6322623E0470180DDB553B10BC422004921548428C41B931081B;
defparam prom_inst_7.INIT_RAM_05 = 256'hB4920371476D26FBBABBA2326F66F66D7FB6B69145008ACB89CF5A0124A3043D;
defparam prom_inst_7.INIT_RAM_06 = 256'hA2F44E8B911A2E5599C76D26DD6671D98842A21A11C3874312C2649869692414;
defparam prom_inst_7.INIT_RAM_07 = 256'h6FF59349BC170DBEF7B5A942F9A228988B07304809249145C9A68A2F44E8BD13;
defparam prom_inst_7.INIT_RAM_08 = 256'h2C60F1C0C1D8CBCC0804504C6E0E0C15526DE5A0415526DE5A041045AAC0CB15;
defparam prom_inst_7.INIT_RAM_09 = 256'h173CDD6749016B0C9DB2693673A010DDF902C9A4DF6AA3860C61334C38BD8810;
defparam prom_inst_7.INIT_RAM_0A = 256'h4B9FDFEF492E7DE8267FC0A9FCBAFB1F35C5146254D532B9E5A3295CD7EC039D;
defparam prom_inst_7.INIT_RAM_0B = 256'h275186349D8AAAAAEECCD249FF7DE5B49A6D4B74B6DAE5F3F3DB6B97DFEFEDD2;
defparam prom_inst_7.INIT_RAM_0C = 256'h9FDCEF3433FE321BA7E73AF91C7C8E2FF46653E7C6EBD73F8EADAFF3F9E799EF;
defparam prom_inst_7.INIT_RAM_0D = 256'h62B47BFBEEFFEC612F33F3EDEFB1097998DD3F39F7E8E3F4717FA3329F3E36AB;
defparam prom_inst_7.INIT_RAM_0E = 256'hCBC92D4102738F274C9834760B142105A5874652439C710F8904F1C71C71C71C;
defparam prom_inst_7.INIT_RAM_0F = 256'hA9D1A80000000000E1F87FFEFFDFBF7FFFFFFFBFFF7FF595823934BEF72F927D;
defparam prom_inst_7.INIT_RAM_10 = 256'h6F5726FF3A64F773F45ECFAB74789B137889896774789B137A800459934D799C;
defparam prom_inst_7.INIT_RAM_11 = 256'hEE72925296B1E00D384E3F2D9B3BCA0E785D59D56F73949294B58F1EAAD9349A;
defparam prom_inst_7.INIT_RAM_12 = 256'h0142A115534CF7D5622B3DF6D642AFCBE49684E336F568CFEF7940CF0B8B3A8D;
defparam prom_inst_7.INIT_RAM_13 = 256'h994BECA5CA6F0EA15AA7BED482C8F4A70D4E5A3087293A529CB5B9C707D02441;
defparam prom_inst_7.INIT_RAM_14 = 256'h2D7DF6FAE0BF0AC14D5F9D2D1DB2DF51D77BB729070084EA6765225220A44A45;
defparam prom_inst_7.INIT_RAM_15 = 256'hA149244A0D6161211425EB8323C370DC143E8770529A12D8EC2612E430C6E415;
defparam prom_inst_7.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0DD423184ED29A0C250;
defparam prom_inst_7.INIT_RAM_17 = 256'h0000FFFFFFFFFFFFFFFF0000FFFFFFFFFFFFFD55FFFEFE9DC2839BFAAC17D06A;
defparam prom_inst_7.INIT_RAM_18 = 256'h00000000000000000000FFFFFFFFFFFF00000FDF000000000400000000000000;
defparam prom_inst_7.INIT_RAM_19 = 256'h0000005144415040A0A6AAAA90561101AAAAAAAAAA9A4403AAAAAAAA712AAAAA;
defparam prom_inst_7.INIT_RAM_1A = 256'h1F5DD74000562503DEB2B242EC76D1E7C749468F9EEF1A9CF8BA5E9202D71FEC;
defparam prom_inst_7.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFAA02A82A08288A208A02A82882A80AA208800;
defparam prom_inst_7.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_7.INIT_RAM_20 = 256'hEBF0052BB07BC7B041044044540001110015004040017FAABF9051AAC12A0782;
defparam prom_inst_7.INIT_RAM_21 = 256'h5541415045144FAFBEE0006BE02B96A541445104540501451504550510545FAF;
defparam prom_inst_7.INIT_RAM_22 = 256'h51441110505550445051000500004FFAEBA0556AA45BD3B44144111450155044;
defparam prom_inst_7.INIT_RAM_23 = 256'hABF0453BA40EC0F451451111505554114004551051410FFAFEA0502AF44E90F0;
defparam prom_inst_7.INIT_RAM_24 = 256'h1551051010040FEFFFB1547BF01ED1E051451111415015110501404545150FFF;
defparam prom_inst_7.INIT_RAM_25 = 256'h50411111054001445054554545405FEEFAA4112BE05A80A45041111101400511;
defparam prom_inst_7.INIT_RAM_26 = 256'hAFC014AEC1EF1EC20411011150000444005401010005FEAAFE4146AB04A81E0A;
defparam prom_inst_7.INIT_RAM_27 = 256'h5505054114513EBEFB8001AF80AE5A9705114411501405145411541441517EBF;
defparam prom_inst_7.INIT_RAM_28 = 256'h45104441415541114144001400013FEBAE8155AA916F4ED30510445140554111;
defparam prom_inst_7.INIT_RAM_29 = 256'hAFC114EE903B03D345144445415550450011544145043FEBFA8140ABD13A43C2;
defparam prom_inst_7.INIT_RAM_2A = 256'h5544144040103FBFFEC551EFC07B478245144445054054441405011514543FFE;
defparam prom_inst_7.INIT_RAM_2B = 256'h41044444150005114151551515017FBBEA9044AF816A02934104444405001444;
defparam prom_inst_7.INIT_RAM_2C = 256'h441043EBEEBD401B50054050105114411405505105501544110003EBFAED554A;
defparam prom_inst_7.INIT_RAM_2D = 256'h1055551450050544115443EABBFD415B50055054105104451415541114144011;
defparam prom_inst_7.INIT_RAM_2E = 256'h54015014145144441055550440411011400557EEBEE9440B5405505414510444;
defparam prom_inst_7.INIT_RAM_2F = 256'h415016FFFEF8511F54015014141144445050054445544005151116EEEBA9444F;
defparam prom_inst_7.INIT_RAM_30 = 256'h4140005110011015040446FFBBAC504F54015014141044445150014115150550;
defparam prom_inst_7.INIT_RAM_31 = 256'h54015014141044444140001050504144515142FBAAEC551B5401501414104444;
defparam prom_inst_7.INIT_RAM_32 = 256'h10410FAFBAF5006E4015014041445104501541441540551044000FAFEBB5552A;
defparam prom_inst_7.INIT_RAM_33 = 256'h415554514014151045510FAAEFF5056F40154150414411145055504450510045;
defparam prom_inst_7.INIT_RAM_34 = 256'h5005405051451110415554110104404500155FBAFBA5102F5015415051441110;
defparam prom_inst_7.INIT_RAM_35 = 256'h05405BFFFBE1447E5005405050451111414015111551001454445BBBAEA5113F;
defparam prom_inst_7.INIT_RAM_36 = 256'h050001444004405410111BFEEEB1413E50054050504111114540050454541541;
defparam prom_inst_7.INIT_RAM_37 = 256'h5005405050411111050000414141051145450BEEABB1546E5005405050411111;
defparam prom_inst_7.INIT_RAM_38 = 256'h0150150150150150150150150150150150140540540540540540540540540540;
defparam prom_inst_7.INIT_RAM_39 = 256'h1501501501501501501501501505405405405405405405405405405405405405;
defparam prom_inst_7.INIT_RAM_3A = 256'h5015015015015015015054054054054054054054054054054054054150150150;
defparam prom_inst_7.INIT_RAM_3B = 256'h0150150150150540540540540540540540540540540540541501501501501501;
defparam prom_inst_7.INIT_RAM_3C = 256'h1501505405405405405405405405405405405405415015015015015015015015;
defparam prom_inst_7.INIT_RAM_3D = 256'hEAFEA54054054054054054054054054050150150150150150150150150150150;
defparam prom_inst_7.INIT_RAM_3E = 256'hAFEAFEAFEAFEAFEAFEAFEAFEAFABFABFABFABFABFABFABFABFABFABFABFABEAF;
defparam prom_inst_7.INIT_RAM_3F = 256'hFEAFEAFEAFEAFEAFEAFABFABFABFABFABFABFABFABFABFABFABFABEAFEAFEAFE;

pROM prom_inst_8 (
    .DO({prom_inst_8_dout_w[30:0],prom_inst_8_dout[4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_8.READ_MODE = 1'b0;
defparam prom_inst_8.BIT_WIDTH = 1;
defparam prom_inst_8.RESET_MODE = "SYNC";
defparam prom_inst_8.INIT_RAM_00 = 256'hFFFFFFFFFFCF3C048834A211A1A22C49FC65E5BFFFFFC59FFEFAFFFFFFFFFF01;
defparam prom_inst_8.INIT_RAM_01 = 256'h8383F16A4C265B1DD7FCEBDCE3F37AA22221FFFF85C813000D0D86F11C210A10;
defparam prom_inst_8.INIT_RAM_02 = 256'hFFFFFFFFFFFA9AB610A50021BAA0A27C934A4B974C3C30010880810284404444;
defparam prom_inst_8.INIT_RAM_03 = 256'h8028C8430165180B2801651142A90ABA124850A1001051400104544110445140;
defparam prom_inst_8.INIT_RAM_04 = 256'h0A94614B30E0A3BDA40D432A80AC04D080014685A5695851A86002128C02528A;
defparam prom_inst_8.INIT_RAM_05 = 256'h4042CC2C2E2E2100B88E1604051010DB16D8808E194150A2128542C4494A14B3;
defparam prom_inst_8.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFC92170820685074684215858444A5142C5452D42C84892909;
defparam prom_inst_8.INIT_RAM_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD49450D142928A093;
defparam prom_inst_8.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_0C = 256'hBBBBBB9B9B0452A569AAA0D5AD56AD6B51102A8A1AB5A8512D456C94AD9AD049;
defparam prom_inst_8.INIT_RAM_0D = 256'hCA81F8CBFB46F3DB64B2C72170D4C907D7131D3C898B04446582262EFDDBBB99;
defparam prom_inst_8.INIT_RAM_0E = 256'h4B636BB4877B7DBB6CA32A07F61B6DB0DB6DF676360A32A07E36CA381F94DB28;
defparam prom_inst_8.INIT_RAM_0F = 256'h1C0A6C02A044830220C0003084934D84870C461202D242BF26856D925124B622;
defparam prom_inst_8.INIT_RAM_10 = 256'hF2FF0FF0F77C3AFB3B318F7B2CDB893499FAB490201B03256DD3B05249641418;
defparam prom_inst_8.INIT_RAM_11 = 256'hA486C920015D699B28932C967094931CB665D45DA124F6773BDDB6CCD44903F2;
defparam prom_inst_8.INIT_RAM_12 = 256'hC0E1620F4EA830130BFEAFFFCE166669B72DCB666F7BDEF7EF7BE38DEF79C35C;
defparam prom_inst_8.INIT_RAM_13 = 256'hDE37045999811862652B3FFA567FF4967FE92CFFD22CFFA42CFF48167E900044;
defparam prom_inst_8.INIT_RAM_14 = 256'h982464AAD320F16666046210002C16666044316666045108000000005858D291;
defparam prom_inst_8.INIT_RAM_15 = 256'h8FC48364FE96DB6C97D73297484B5E9BB2492DBB9098E2E5F5B158899DDB9599;
defparam prom_inst_8.INIT_RAM_16 = 256'hFFFFFFC0A5790EFFFFBFC8F0307BBBF2EEFCBF7E4AFE57E6DCD3B65DF53EA1BD;
defparam prom_inst_8.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_8.INIT_RAM_18 = 256'hA02A0280A028282820A28A2882222222208282A000282220008A0000755FD77C;
defparam prom_inst_8.INIT_RAM_19 = 256'h0C4AAAAAA800002AAAA0000AAAA0002AAA000AAA000AA800AA802A802A80AA02;
defparam prom_inst_8.INIT_RAM_1A = 256'hF920E9312548BB6000749F0A5E78520D2EB4922A9202D2A42BA020000C482000;
defparam prom_inst_8.INIT_RAM_1B = 256'hDB74CDC07DADC04EB6DC1249C6D72BEDAE095B111E178737094A8FCB55AA07EA;
defparam prom_inst_8.INIT_RAM_1C = 256'h00811B321032EF2C3A34B20C6CD9C4096312D92649D6B373499B094D0C9B3007;
defparam prom_inst_8.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF4F49A736C9EB;
defparam prom_inst_8.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_8.INIT_RAM_20 = 256'hDFF37FDFF9357EFFF9ABF7FF357BFF9ABDFF357B63BAF5111B97000454110440;
defparam prom_inst_8.INIT_RAM_21 = 256'hDAE6E9592AC9544AB255929F4250CA7420B4BDFFCDFF7FF9357BFE6FFEFFC9AB;
defparam prom_inst_8.INIT_RAM_22 = 256'h8981845C84C11C814514AA0F251052883C8D6D6E6DC0AA21441E0A20A550791A;
defparam prom_inst_8.INIT_RAM_23 = 256'h44C086DE44C20E470D70C12811302DA393309BC8C1C2504D348239334D1C8C9A;
defparam prom_inst_8.INIT_RAM_24 = 256'h330889BC8C1C25489A3690464721364D11C8809934218820A4441C8C49191C88;
defparam prom_inst_8.INIT_RAM_25 = 256'h74F3D26D3CF4F080242126690C2226F2330888391C35C304A80826610D134472;
defparam prom_inst_8.INIT_RAM_26 = 256'h7499D2731D3C674B1B4F19D3C2009482010406D274F3D371D2F4F134F3D2F4DC;
defparam prom_inst_8.INIT_RAM_27 = 256'hB56945142A8F055042A83C8D6D7369E00411313491D3CC74DC67499D3CE4D3C6;
defparam prom_inst_8.INIT_RAM_28 = 256'hA03D276CF7A789A7B7410009A7B67BD271D3DB8114508A3C14414AA0F235B5CD;
defparam prom_inst_8.INIT_RAM_29 = 256'h7B7082011134F6CF33A6E33A7B70210F4F6C7369E7A7ADD09E9EB63BD3C749DB;
defparam prom_inst_8.INIT_RAM_2A = 256'h67A0084023A7B679134F39D3D6E8CE9EB6799D3CC749DBA111D376C733A79C9A;
defparam prom_inst_8.INIT_RAM_2B = 256'h9E04749C74F6E0E9ED8ECD3DBA769ED9E8221334F3D3C6E9E9EB639D3DB83A7B;
defparam prom_inst_8.INIT_RAM_2C = 256'h8074F1D376E0E9BB67BD3D6E9E9E363810053D3CED3DB8669ED8EF4DDB87A4ED;
defparam prom_inst_8.INIT_RAM_2D = 256'hDD31D3DB3CCDA7B7466D3DB1D20880C4D3C474F1BA23A78D9EE74F6E9CE9ED8E;
defparam prom_inst_8.INIT_RAM_2E = 256'hEB70E74F1B3C0900519D3CE6D3DB87369ED8EC749DB873A4ED9E0488E9B98E9E;
defparam prom_inst_8.INIT_RAM_2F = 256'hDA1D499C4C3AFBACD8D4DDD606E35A5E77BA3D09263A78CE93B706749DB3DCE9;
defparam prom_inst_8.INIT_RAM_30 = 256'h5656DAD67A1E8F4743D8F63D8F69F4D9C69D7DD66BA6EE1B1E87A3D2E93D8F63;
defparam prom_inst_8.INIT_RAM_31 = 256'hEB33A4B3F67D9DAE97E8FA3D1D24B5371E759B3DBA771AD4DC79D66CE9D6A35A;
defparam prom_inst_8.INIT_RAM_32 = 256'h75F732D276F533AFB99695A8F7ECFB3D9D9FA3E8F474D749C79D64D338FA6EBE;
defparam prom_inst_8.INIT_RAM_33 = 256'h0F43D0F47492D49C775DB56A4EBBAC8E974EB1E87A1E87A5D27B1EC7B1EDD6A6;
defparam prom_inst_8.INIT_RAM_34 = 256'h43D2E93D8F63D8F63DB2D4DC71E7592725A938E3CEB24D6A3CF63D8F69ECED3D;
defparam prom_inst_8.INIT_RAM_35 = 256'h9ECED74BA496A6EB8F3AC99216A4E38FBB75921E87A1E87A1E8E9D63D0F43D0F;
defparam prom_inst_8.INIT_RAM_36 = 256'hF4BA4F6CB5375C79D3AC9392D49C71F76EB363D8F63D8F63DB7B8F3D8F63D8F6;
defparam prom_inst_8.INIT_RAM_37 = 256'h92D4DD75F74EB36485A938EBEEDD66EC7A1E87A1E87A1E8E9D63D0F43D0F43D0;
defparam prom_inst_8.INIT_RAM_38 = 256'hB759B2725A938EBEEDD66EC7B1EC7B1EC7B1EDBDC79EC7B1EC7B1ED3D9DAE974;
defparam prom_inst_8.INIT_RAM_39 = 256'hD77DD3ACD90F43D0F43D0F43D0F474CB1E87A1E87A1E87A1E9749ED96A6EBAFB;
defparam prom_inst_8.INIT_RAM_3A = 256'hF63D8F63D8F69EA3CF63D8F63D8F63DA7B3B5D2E9A7A938E3BEEDD66ED8F5275;
defparam prom_inst_8.INIT_RAM_3B = 256'hD0F43D0F43D0F43D0F4BA4F6EF5271C77DDBACDDBDBD49D75DE74EB2738F63D8;
defparam prom_inst_8.INIT_RAM_3C = 256'h97492D4DC719E776EB376C5A9BAEBBCCE9D64C87A1E87A1E87A1E87A1E8E9D63;
defparam prom_inst_8.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9EC7B1EC7B1EC7B1ED3D9DAE;
defparam prom_inst_8.INIT_RAM_3E = 256'h0000FFFFFF000000FFFFFF000000FFFFFF000000FFFFFF000000FFFFFF000000;
defparam prom_inst_8.INIT_RAM_3F = 256'hFFFFFF000000FFFFFF000000FFFFFF000000FFFFFF000000FFFFFF000000FFFF;

pROM prom_inst_9 (
    .DO({prom_inst_9_dout_w[30:0],prom_inst_9_dout[4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_9.READ_MODE = 1'b0;
defparam prom_inst_9.BIT_WIDTH = 1;
defparam prom_inst_9.RESET_MODE = "SYNC";
defparam prom_inst_9.INIT_RAM_00 = 256'h0C34D34D35822CD24A5B608B445440192918760855EA862C128000410000012D;
defparam prom_inst_9.INIT_RAM_01 = 256'h1252481999E66679999E66663EEEF6FFE6660F8EEF6FFE6620EB664289441041;
defparam prom_inst_9.INIT_RAM_02 = 256'h25B4D34CB6906C69A5B5A360DDF65461CA95080DA2C2C8BBBB999999F9DFE3F0;
defparam prom_inst_9.INIT_RAM_03 = 256'hCD02ADC590246646AA63676C55663676C55663676C556F12095552F120955525;
defparam prom_inst_9.INIT_RAM_04 = 256'h8904AAA91548C7496AB49565619F07771920CCCAE496DB676B5B9E54BB2B2832;
defparam prom_inst_9.INIT_RAM_05 = 256'hA924076569F8FC7FFEEEEEFFDB7DB7DB616DB55741BADBD92A24536DA6824977;
defparam prom_inst_9.INIT_RAM_06 = 256'hA0DD5E83757A0DD585D5F8FC7D617578904AAA9154971A4790D4ECD948524804;
defparam prom_inst_9.INIT_RAM_07 = 256'hD964FE3F148B2D90852908D269922159D3365148475D7541BA69AA0DD5E83757;
defparam prom_inst_9.INIT_RAM_08 = 256'h2149039595A2BA98585245CC0CACAC333FE5E584C333FE5E584C71C7E2C4890C;
defparam prom_inst_9.INIT_RAM_09 = 256'hB05ACD6892008F080FEFC7E34B811295D122BF1F85F828234545766CA59CA112;
defparam prom_inst_9.INIT_RAM_0A = 256'hDA62E5CB5B699B6965DB88A5FBA0D93E818C1462509422B5E512E939CF242359;
defparam prom_inst_9.INIT_RAM_0B = 256'hC3A388748CBB99BBFFDDFFFFAA6DBFBFF7FF4DB7F5B69ABD7AD6DA6AE5CB3DB6;
defparam prom_inst_9.INIT_RAM_0C = 256'h8F43393F0CE2686BDB2620193C8D9F2A14F6D3E3EEDBB71E894651F0FC772EF2;
defparam prom_inst_9.INIT_RAM_0D = 256'h46140BCA0400408504C3C204108228264B5ED83120E9E47CF940A7B69F1F7423;
defparam prom_inst_9.INIT_RAM_0E = 256'h89C510A914ABA424A9B242E23A1ACC51D5B46CEADB5D222CD388E18618618618;
defparam prom_inst_9.INIT_RAM_0F = 256'h1881840000000000735CD554AA952A555555552AAA544C1525B7EAD062008A18;
defparam prom_inst_9.INIT_RAM_10 = 256'hDBE4FC60953FD910EB686B652FE7F4FF2B699DAD2FE7F4FF2B681B6B7E2C01D1;
defparam prom_inst_9.INIT_RAM_11 = 256'hCC421FC85005563A65E971FC0D0F4F08F2477D57666210FE42802AA599CFE3F1;
defparam prom_inst_9.INIT_RAM_12 = 256'h966A452510205FF5464E17FDB5E3A02B92F15E9713F56E3E35E9E01E48CFAACC;
defparam prom_inst_9.INIT_RAM_13 = 256'h4D714EBBEBAF44ED3282FF95818ECBEE0485DEE29EF7F5CFB81214B222848485;
defparam prom_inst_9.INIT_RAM_14 = 256'hAE4BA0D59B95C1008C0AC8064A1B9939257AB240BE187EA88FB5D35D3ABA6BA7;
defparam prom_inst_9.INIT_RAM_15 = 256'hEA7DB6055F030303268D7AB901E0F81E0D37B67834BED5B8DC2E36FD35C04465;
defparam prom_inst_9.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBDF9E6318DCF7D55C672;
defparam prom_inst_9.INIT_RAM_17 = 256'h000000000000000000000000FFFFFFFF00000D8E000002421E19E00CC94FE526;
defparam prom_inst_9.INIT_RAM_18 = 256'h0000000000000000000000000000000000000C00000000000000000000000000;
defparam prom_inst_9.INIT_RAM_19 = 256'hFFFFFFABFAFBEBBF0E0800003EF8EAAB000000000030AEA8000000008FC00000;
defparam prom_inst_9.INIT_RAM_1A = 256'h2088001F5DD2A3038F42AA60CE2594F34248D5873A4C541E689DF924011E1B76;
defparam prom_inst_9.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFAA0002AA02A82A08288A208A02A82882A80AA;
defparam prom_inst_9.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_9.INIT_RAM_20 = 256'h555FAFEBF0052BB115014141444444140001110011004040417FAABF9051AAD1;
defparam prom_inst_9.INIT_RAM_21 = 256'h5540445541415045144FAFBEE0006BE015415041444144501501440504541510;
defparam prom_inst_9.INIT_RAM_22 = 256'h05415051441114505550445051000540000FFAEBA0556AA01541505144511450;
defparam prom_inst_9.INIT_RAM_23 = 256'h150FFFAAF0453AA405405050441110415554114004551015410FFAFEA0502AF4;
defparam prom_inst_9.INIT_RAM_24 = 256'h4005141551041010154EEFFFF4507BF005405050451111415055110541404545;
defparam prom_inst_9.INIT_RAM_25 = 256'h05405050411111050001445014554545405FEEFAA4112BE00540505045111141;
defparam prom_inst_9.INIT_RAM_26 = 256'h557EBFAFC014AEC55405050511111050000444004401010105FEAAFE4146AB44;
defparam prom_inst_9.INIT_RAM_27 = 256'h5501115505054114513EBEFB8001AF8055054105110511405405101411505441;
defparam prom_inst_9.INIT_RAM_28 = 256'h15054145104451415541114144001500003FEBAE8155AA815505414511445141;
defparam prom_inst_9.INIT_RAM_29 = 256'h543FFEABC114EA9015014141104441055550450011544055043FEBFA8140ABD1;
defparam prom_inst_9.INIT_RAM_2A = 256'h0014505544104040553BBFFFD141EFC015014141144445054154441505011514;
defparam prom_inst_9.INIT_RAM_2B = 256'h15014141044444140005114051551515017FBBEA9044AF811501414114444505;
defparam prom_inst_9.INIT_RAM_2C = 256'h144011441043EBEE50001550055054105114411405505105501544114003EBFA;
defparam prom_inst_9.INIT_RAM_2D = 256'h5144441055551450051544115443EABB50000554055054145104451415541114;
defparam prom_inst_9.INIT_RAM_2E = 256'h54000554015014145144441055150441411011400557EEBE5400055401505414;
defparam prom_inst_9.INIT_RAM_2F = 256'h151550515016FFFE54000554015014141144445050014445544105151117EEEB;
defparam prom_inst_9.INIT_RAM_30 = 256'h1044444140005110011015040446FFBB54000554015014141044445140004115;
defparam prom_inst_9.INIT_RAM_31 = 256'h54000554015014141044444100501050504144515146FAAA5400055401501414;
defparam prom_inst_9.INIT_RAM_32 = 256'h51004510410FAFBA4000554015415041445104501541441540551045000FAFEB;
defparam prom_inst_9.INIT_RAM_33 = 256'h451110415554514014551045510FAAEE40001550154150514411145055504450;
defparam prom_inst_9.INIT_RAM_34 = 256'h5000155005405051451110415454110504404500155FBAFB5000155005415051;
defparam prom_inst_9.INIT_RAM_35 = 256'h54554145405BFFFB5000155005405050451111414005111551041454445FBBAE;
defparam prom_inst_9.INIT_RAM_36 = 256'h411111050001444004405410111BFEEE50001550054050504111114500010454;
defparam prom_inst_9.INIT_RAM_37 = 256'h5000155005405050411111040140414141051145451BEAAB5000155005405050;
defparam prom_inst_9.INIT_RAM_38 = 256'h5400155400155400155400155400155400155000555000555000555000555000;
defparam prom_inst_9.INIT_RAM_39 = 256'h4001554001554001554001554005550005550005550005550005550005550005;
defparam prom_inst_9.INIT_RAM_3A = 256'h0015540015540015540055500055500055500055500055500055500155400155;
defparam prom_inst_9.INIT_RAM_3B = 256'h0155400155400555000555000555000555000555000555001554001554001554;
defparam prom_inst_9.INIT_RAM_3C = 256'h1554005550005550005550005550005550005550015540015540015540015540;
defparam prom_inst_9.INIT_RAM_3D = 256'h5500055500055500055500055500055500155400155400155400155400155400;
defparam prom_inst_9.INIT_RAM_3E = 256'h5000555000555000555000555001554001554001554001554001554001554005;
defparam prom_inst_9.INIT_RAM_3F = 256'h0005550005550005550015540015540015540015540015540015540055500055;

pROM prom_inst_10 (
    .DO({prom_inst_10_dout_w[30:0],prom_inst_10_dout[5]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_10.READ_MODE = 1'b0;
defparam prom_inst_10.BIT_WIDTH = 1;
defparam prom_inst_10.RESET_MODE = "SYNC";
defparam prom_inst_10.INIT_RAM_00 = 256'hFFFFFFFFFFDFFFFDFBFFFEFBFFD1FFFEFD60E0FFFFFFA4A000FEFFFFFFFFFFC1;
defparam prom_inst_10.INIT_RAM_01 = 256'hC58FF1E88EE4C30FDBBCC64EC4E23FA051FA00008408C9FFFFFEFDFFFE1FFDFE;
defparam prom_inst_10.INIT_RAM_02 = 256'hFFFFFFFFFFFE19934F86EFF43B88C87473CE088A0C002FF1223FFFFFFD51FFFF;
defparam prom_inst_10.INIT_RAM_03 = 256'h8402E9C572605B9302426044100440189B6D4408555541555405105444051405;
defparam prom_inst_10.INIT_RAM_04 = 256'hA0917448BA5A038892A4100A4A2EA1C1D024169FA3E8FD05F8AE42702DCA302F;
defparam prom_inst_10.INIT_RAM_05 = 256'h1080258585858A02012C1C1C8344A409C04E212D74CCDA1A3820106168C0859B;
defparam prom_inst_10.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFF418825234C29470C00081A0F174704101011381069E2D1D18;
defparam prom_inst_10.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF09C73F1CE138E412;
defparam prom_inst_10.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_0C = 256'h99BBBB9B9800C28624922945AC4A2D621C5578E248B5809564716D90A8024809;
defparam prom_inst_10.INIT_RAM_0D = 256'h820E4A2496D0B6D240644305604847F3B60855992AAB495D5DA4AEAF4FF9D9BB;
defparam prom_inst_10.INIT_RAM_0E = 256'hC81027F685004D1A4822083934124920924934B4F402208393248220E4849208;
defparam prom_inst_10.INIT_RAM_0F = 256'h582A6E6BF4666B530AE8FF8890C2CC0CBEA4D2B100032B9104572083146588AA;
defparam prom_inst_10.INIT_RAM_10 = 256'hC3DB15B153EE615F5EA10C701DFF0190C8DA6D10927F068726C990C32522B248;
defparam prom_inst_10.INIT_RAM_11 = 256'h95A25B72594D64A965B96DB2E9BDB74D932CC84CA107C40743A1B6C4105BAFF7;
defparam prom_inst_10.INIT_RAM_12 = 256'hC9A1CC5E9DCC1D9909B6A8C0041E6669360D83666C6318C60C63030D8C6083FC;
defparam prom_inst_10.INIT_RAM_13 = 256'h226085CCCCC699D042894001128002128004250008250010250020128040004C;
defparam prom_inst_10.INIT_RAM_14 = 256'hCC701D95BDA4F733331A6437FF01733331A4B733331A5213FFFFFFFE06793E6B;
defparam prom_inst_10.INIT_RAM_15 = 256'h1A4406C4DA96DB6DB7172375B6DC1A18968B6FB3588000007000007EEAA984CC;
defparam prom_inst_10.INIT_RAM_16 = 256'hFFFFFF8086658A0000401304C44200848021081093FE5786D852B6BDFF7CCB3E;
defparam prom_inst_10.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_10.INIT_RAM_18 = 256'hA000AA800AA802A80AA02A0280A0A0A0A28A2088888A282AAA8200000A082080;
defparam prom_inst_10.INIT_RAM_19 = 256'h1180AAAAA8000000000AAAAAAAA0000000AAAAAA000002AAAA80002AAA8000AA;
defparam prom_inst_10.INIT_RAM_1A = 256'h24FE4430892AD96C194C47A11668C9656594566031004320A93E0C0011800C00;
defparam prom_inst_10.INIT_RAM_1B = 256'h28C3531F82934E91A49180970598042310C09880012840245208B404880FF813;
defparam prom_inst_10.INIT_RAM_1C = 256'h0DF2BB35309072CD564C85CC6CD98BF2D4A2496C5B34D000D206D208BC0641F8;
defparam prom_inst_10.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF46022436DB8B;
defparam prom_inst_10.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_10.INIT_RAM_20 = 256'h02040801024300040218008043001021802043003CC603FE33B0000EBAEAAFAE;
defparam prom_inst_10.INIT_RAM_21 = 256'hBE75DC984482261130890402F08C0413FCBD8008102001024300408040081218;
defparam prom_inst_10.INIT_RAM_22 = 256'h220F1DA1D10761D2773D339B4D98E4EC6DED5F272BA6EC7277369BB9C99CDBDA;
defparam prom_inst_10.INIT_RAM_23 = 256'h990F1D30E50EF0E70770C1383443CA6C3943E61CC1C27D194E0EC3967361CC8F;
defparam prom_inst_10.INIT_RAM_24 = 256'h6633B261CC1C27F232C9C19F98746793E61D81D91F5A20CF39F9E1D10E7661C8;
defparam prom_inst_10.INIT_RAM_25 = 256'h0C843393210C80802623E88679CFD9874433B3C39C1DC304FC1F6CCE71ECF987;
defparam prom_inst_10.INIT_RAM_26 = 256'h8CC63386E32138CC64C8463202009C82010499330C863384330C844C84330CE1;
defparam prom_inst_10.INIT_RAM_27 = 256'hAF5A763DB39B4D98F4CC6DED5F395C380412464CEE32138CE1B8CE63211B321B;
defparam prom_inst_10.INIT_RAM_28 = 256'h2343280788642664004101226403C4338432004D98E4EE6DA7739339B7B57CE5;
defparam prom_inst_10.INIT_RAM_29 = 256'h400C8202464C8078DC6709C640002198C80788990C643011A19043863218CE00;
defparam prom_inst_10.INIT_RAM_2A = 256'h38200874CC640384ECC86E32081B3190C386E32118CE00226E328070CC642366;
defparam prom_inst_10.INIT_RAM_2B = 256'hE00D8CA18C801B1900E1932006C9900E0822364C86321813190C384320068640;
defparam prom_inst_10.INIT_RAM_2C = 256'h898C8632801B19C038632081B190C3C010076321932006D9900E18CA006C6700;
defparam prom_inst_10.INIT_RAM_2D = 256'h026E3201E27664009193201C3208891932138C86068C6410E118C801A71900F0;
defparam prom_inst_10.INIT_RAM_2E = 256'h040998C861E0110074632119320069D9900E138CA0069C6700E0093319433190;
defparam prom_inst_10.INIT_RAM_2F = 256'hB9A2CA209D813439A72CA209DACB56D9632D011A4CC643319C00998CA01E3719;
defparam prom_inst_10.INIT_RAM_30 = 256'hD966BC64160582C2C0B82E0B82E98CA20C809A1CD86510C9058160B0580B82E0;
defparam prom_inst_10.INIT_RAM_31 = 256'h0E7964902E0B8B858058160B0B33CB282787348B9218272CE19E1CF658D2CB56;
defparam prom_inst_10.INIT_RAM_32 = 256'h8268613309CB3C13430993B4005C170B8B8160582C2CD8CA09A1CD90C3C6504D;
defparam prom_inst_10.INIT_RAM_33 = 256'h02C0B02C2C8F2CE1882277167044136582C4905816058160B01705C1705CD967;
defparam prom_inst_10.INIT_RAM_34 = 256'hC0B0580B82E0B82E0B922CE1867873D8DC59C30CF0E7BDAD002E0B82E05C5C0B;
defparam prom_inst_10.INIT_RAM_35 = 256'h05C5C2C16639650413439A2779650413C38734858160581605858920B02C0B02;
defparam prom_inst_10.INIT_RAM_36 = 256'h2C1602E6CB28209A1439A4272CA0827870E7B0B82E0B82E0BA4B400B82E0B82E;
defparam prom_inst_10.INIT_RAM_37 = 256'h862CA0826850E6899C59410CF0E1CF3616058160581605858DA0B02C0B02C0B0;
defparam prom_inst_10.INIT_RAM_38 = 256'h28734484E59410CF0E1CF361705C1705C1705D25A005C1705C1705C0B8B8582C;
defparam prom_inst_10.INIT_RAM_39 = 256'h199E1C39E6C2C0B02C0B02C0B02C2C490581605816058160582C05CD96504134;
defparam prom_inst_10.INIT_RAM_3A = 256'h2E0B82E0B82E929002E0B82E0B82E0B817170B0590C59C30C4D0A1CD1338B286;
defparam prom_inst_10.INIT_RAM_3B = 256'hB02C0B02C0B02C0B02C1602E48B386189A1439A24262CA18667870E79902E0B8;
defparam prom_inst_10.INIT_RAM_3C = 256'h82CC72CE186678850E689DE59C30CCF30E1CF3616058160581605816058589A0;
defparam prom_inst_10.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF85C1705C1705C1705C0B8B85;
defparam prom_inst_10.INIT_RAM_3E = 256'hFFFF000000000000FFFFFFFFFFFF000000000000FFFFFFFFFFFF000000000000;
defparam prom_inst_10.INIT_RAM_3F = 256'hFFFFFFFFFFFF000000000000FFFFFFFFFFFF000000000000FFFFFFFFFFFF0000;

pROM prom_inst_11 (
    .DO({prom_inst_11_dout_w[30:0],prom_inst_11_dout[5]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_11.READ_MODE = 1'b0;
defparam prom_inst_11.BIT_WIDTH = 1;
defparam prom_inst_11.RESET_MODE = "SYNC";
defparam prom_inst_11.INIT_RAM_00 = 256'h6DB6DB6DB70A2656DACBE01F09F0092FBC06BE0100FFD76A137FFFC6FFFF0921;
defparam prom_inst_11.INIT_RAM_01 = 256'h809B25BBB9AEEF6BBBDAEEE66276FEEEEE661C876FEEEEE72BCFE6019B2DB6DB;
defparam prom_inst_11.INIT_RAM_02 = 256'h2000410E11B62220808DB114C46702AA5645A3418A6888BBBBBBBB99D9FB7DBE;
defparam prom_inst_11.INIT_RAM_03 = 256'h4D0004C48912152C00312364C02312364C02312364C029101B54069101B54060;
defparam prom_inst_11.INIT_RAM_04 = 256'h880DAA033018C74520144020319D29331901ADDA6DB2493329499E4089096210;
defparam prom_inst_11.INIT_RAM_05 = 256'h300019E025F8FC5776666676D92D92D9206D93D0E89848CA0169412492662034;
defparam prom_inst_11.INIT_RAM_06 = 256'hF44C07D1301F44C5A481F8FC31E9204880DAA03301831AE79442244B1E60002F;
defparam prom_inst_11.INIT_RAM_07 = 256'hFBECB61B120F1F90842948C6798E605B83870402030C30E898618744C07D1301;
defparam prom_inst_11.INIT_RAM_08 = 256'h6801A38080902088080A20E48404043336E5F5ADC3336E5B7ADC30C36AC199CC;
defparam prom_inst_11.INIT_RAM_09 = 256'h901521E0000053A50B66C36082A8300553079B0D80DB710A1000122581CCB037;
defparam prom_inst_11.INIT_RAM_0A = 256'hDE22C58BDB78993BED4A81E5BBE04FBE00873D26BDAF69757B76E7CBDB6406CB;
defparam prom_inst_11.INIT_RAM_0B = 256'hD564CC7F8C99999DDDFFF6DB22CFF6FDBEDBDB249DB788B162F6DE22C58B6FB6;
defparam prom_inst_11.INIT_RAM_0C = 256'hAE31066C845CE0713122631222081013108E0B4B5C48975C085810A4522B072C;
defparam prom_inst_11.INIT_RAM_0D = 256'h566D2B420EC46AA778434A0D88AA3BC20B8989133AB11150809A84705A5AE403;
defparam prom_inst_11.INIT_RAM_0E = 256'hC79441E94A79EC356C306BE20236ED45D5B4227A5ACB6364D15A410410410410;
defparam prom_inst_11.INIT_RAM_0F = 256'h5CC49400000000000A42911222448904104104820904B2FD86B369B5FF1021FF;
defparam prom_inst_11.INIT_RAM_10 = 256'hFD546C05142DB772B6DC1FED3CC1B53732C7D3613CC1B53732CE56D8361883C1;
defparam prom_inst_11.INIT_RAM_11 = 256'hAAABBBFEFDAFB00921E9F427DD694825E8A51B1D4D555DDFF7ED7D87BBCB61B0;
defparam prom_inst_11.INIT_RAM_12 = 256'hE22FCD7538B84DB54EE6136FF552A07DD7F51E9F15B548A7752905BD14A363A9;
defparam prom_inst_11.INIT_RAM_13 = 256'h48515C2AC2B7046C92426DD2808C6BFF4505C8E6BEEFECCFFD1410A26A427ED4;
defparam prom_inst_11.INIT_RAM_14 = 256'h66112D93A04414A4EC8A89650997591525DEFA29770ABDBAB3215615682AC2AC;
defparam prom_inst_11.INIT_RAM_15 = 256'h242FFFC00C14141561B7FFB314F43D2F44FE9F7D119A321D0EC751F4F4EFE134;
defparam prom_inst_11.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF790014A50856C00EA10;
defparam prom_inst_11.INIT_RAM_17 = 256'h0000FFFFFFFFFFFFFFFF000000000000FFFFF218FFFFFF7A642CABFD5B3FF9B4;
defparam prom_inst_11.INIT_RAM_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_11.INIT_RAM_19 = 256'h5555554100010145555155555541415455555555455505555555555541555555;
defparam prom_inst_11.INIT_RAM_1A = 256'h2A80AA20880353CBAEFE66AACAA59AEBF36EE9D75F6DA75D7E04480000A75D11;
defparam prom_inst_11.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF80AAAAAA0002AA02A82A08288A208A02A8288;
defparam prom_inst_11.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_11.INIT_RAM_20 = 256'h551510555FAFEBF000554015414141044444140005110011004040417FAABF90;
defparam prom_inst_11.INIT_RAM_21 = 256'h1104505540445541415045144FAFBEE000155015414041445144500501451504;
defparam prom_inst_11.INIT_RAM_22 = 256'h00155005415051441114505550445011004540000FFAEBA00015500541505144;
defparam prom_inst_11.INIT_RAM_23 = 256'h404545150FFFABF000155005415051451110415554114004551015410FFAFEA0;
defparam prom_inst_11.INIT_RAM_24 = 256'h1111454005151551151010150FEFFFF400155005405050451111415015110541;
defparam prom_inst_11.INIT_RAM_25 = 256'h00155005405050411111050001445014554545405FEEFAA40015500540505045;
defparam prom_inst_11.INIT_RAM_26 = 256'h545441557EBFAFC00155005505050411111050001444004401010105FEAAFE41;
defparam prom_inst_11.INIT_RAM_27 = 256'h4411415501115505054114513EBEFB8000554055050105114511401405145411;
defparam prom_inst_11.INIT_RAM_28 = 256'h00554015054145104451415541114044011500003FEBAE810055401505414510;
defparam prom_inst_11.INIT_RAM_29 = 256'h011514543FFEAFC100554015054145144441055550450011544055043FEBFA81;
defparam prom_inst_11.INIT_RAM_2A = 256'h4445150014545544544040543FBFFFD100554015014141144445054054441505;
defparam prom_inst_11.INIT_RAM_2B = 256'h00554015014141044444140005114051551515017FBBEA900055401501414114;
defparam prom_inst_11.INIT_RAM_2C = 256'h5411141440114410055555500005540550541051144114055051055055441140;
defparam prom_inst_11.INIT_RAM_2D = 256'h5014145144441055550450051544115405555554000554015054145104451415;
defparam prom_inst_11.INIT_RAM_2E = 256'h0155555400055401501414514444105415044141101140050155555400055401;
defparam prom_inst_11.INIT_RAM_2F = 256'h0051150515505150015555540005540150141411444450500145455441041511;
defparam prom_inst_11.INIT_RAM_30 = 256'h5014141044444140005110011015040401555554000554015014141044445140;
defparam prom_inst_11.INIT_RAM_31 = 256'h0155555400055401501414104414410050105050414051510155555400055401;
defparam prom_inst_11.INIT_RAM_32 = 256'h5044505100451041155555400015501541504144510450154144154155104500;
defparam prom_inst_11.INIT_RAM_33 = 256'h4050514511104155541140145510455115555550001550054150514411145055;
defparam prom_inst_11.INIT_RAM_34 = 256'h0555555000155005405051451110415054110504404500150555555000155005;
defparam prom_inst_11.INIT_RAM_35 = 256'h0144541455414540055555500015500540505045111141400515155104105444;
defparam prom_inst_11.INIT_RAM_36 = 256'h4050504111110500014440044054101105555550001550054050504111114500;
defparam prom_inst_11.INIT_RAM_37 = 256'h0555555000155005405050411051040140414141050145450555555000155005;
defparam prom_inst_11.INIT_RAM_38 = 256'h0000155555400000155555400000155555400000555555000000555555000000;
defparam prom_inst_11.INIT_RAM_39 = 256'h5554000001555554000001555550000005555550000005555550000005555550;
defparam prom_inst_11.INIT_RAM_3A = 256'h0015555540000015555500000055555500000055555500000055555400000155;
defparam prom_inst_11.INIT_RAM_3B = 256'h5400000155555000000555555000000555555000000555554000001555554000;
defparam prom_inst_11.INIT_RAM_3C = 256'h1555550000005555550000005555550000005555540000015555540000015555;
defparam prom_inst_11.INIT_RAM_3D = 256'h0000055555500000055555500000055555400000155555400000155555400000;
defparam prom_inst_11.INIT_RAM_3E = 256'h5555000000555555000000555554000001555554000001555554000001555550;
defparam prom_inst_11.INIT_RAM_3F = 256'h0005555550000005555540000015555540000015555540000015555500000055;

pROM prom_inst_12 (
    .DO({prom_inst_12_dout_w[30:0],prom_inst_12_dout[6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_12.READ_MODE = 1'b0;
defparam prom_inst_12.BIT_WIDTH = 1;
defparam prom_inst_12.RESET_MODE = "SYNC";
defparam prom_inst_12.INIT_RAM_00 = 256'hFFFFFFFFFFC000FEFC76FF3C0FEEFF6FFDC5C5FFFFFFBD801EF9FFFFFFFFFF87;
defparam prom_inst_12.INIT_RAM_01 = 256'h8319A3238420144DAF746A58C3D17189339255551100D300107FFE01FFE33E7F;
defparam prom_inst_12.INIT_RAM_02 = 256'hFFFFFFFFFFFEB3965EB16BB198AE3F20C92062D365B5AFF10440810204624444;
defparam prom_inst_12.INIT_RAM_03 = 256'hD4ABE56F3B7579DBABEB75755AA96AA2F6DC16AD554501555550110005054005;
defparam prom_inst_12.INIT_RAM_04 = 256'h2A56653B32D2A129B23D592AC89932C8C8355E5595655C57DDE7491ABCE91ABD;
defparam prom_inst_12.INIT_RAM_05 = 256'h5B58A42424242D64A1B6C6C53196D60B105899B75D5544B95AB55AF5E46AD2A3;
defparam prom_inst_12.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFEC2D77B82EBF722E96AD63595C2B565A995C8D5AE46BC8C8D;
defparam prom_inst_12.INIT_RAM_07 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_12.INIT_RAM_08 = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_12.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF64D37B4DEC9A6EC9;
defparam prom_inst_12.INIT_RAM_0A = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_12.INIT_RAM_0B = 256'h5555555555555555555555555555555555555555555555555555555555555555;
defparam prom_inst_12.INIT_RAM_0C = 256'hCC888888888A59B1DA456CD7BD66BDEB5179A2893AF7A408A1459C4632A52164;
defparam prom_inst_12.INIT_RAM_0D = 256'h954ADE7DB6F2B0DB78338C20312527389012004C999864C4C43262628CCC8888;
defparam prom_inst_12.INIT_RAM_0E = 256'h5A8D92185D086D9B6D5A552B72DB6DB6DB6D86060655A552B7B6D5A4ADAADB56;
defparam prom_inst_12.INIT_RAM_0F = 256'hE38D3316B72E0CB703362AD6660BFEE5867A694AA218404CB080875838AC2833;
defparam prom_inst_12.INIT_RAM_10 = 256'hDADBEDBEDB6D6CDB3E2D6DFCEC5B6C462EDD6F55DD0B92D8D8366258DA9C6DF1;
defparam prom_inst_12.INIT_RAM_11 = 256'hCB1DB6C010341B161B66D30C27670C306CC331622BB0D8B3198CB6D22ADB85B0;
defparam prom_inst_12.INIT_RAM_12 = 256'hF5C1F6C95DFC408EDD9718C05A072333966599622C6318C60C6309258C6B411D;
defparam prom_inst_12.INIT_RAM_13 = 256'h328AB3D999F2BCFB16FB0079F600F3F601E7EC03CF6C079E6C0F3C361E7800C1;
defparam prom_inst_12.INIT_RAM_14 = 256'h9F118C6C77325F6667CAF3C155D8F6667CA21F6667CAC9E8AAAAAAABB2CE19BC;
defparam prom_inst_12.INIT_RAM_15 = 256'h7E6D13DDCBB6DB6DB66666C3ECDE4ECDB75B70CC9E528A8D25A55288888B1D99;
defparam prom_inst_12.INIT_RAM_16 = 256'hFFFFFFFDB029E10000000C03030240849021081092663BB6DB765215BCEDF82D;
defparam prom_inst_12.INIT_RAM_17 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_18 = 256'h0AAAAA800002AAA8000AAA002AA00AA00A80A0282828A20888A2000020288801;
defparam prom_inst_12.INIT_RAM_19 = 256'h0E7EAAAAA800000000000000000AAAAAAAAAAAAA00000000002AAAAAAA800000;
defparam prom_inst_12.INIT_RAM_1A = 256'h90E72D96E44004B1E01A532B722E7658186FA98ACAA25804040622800E7C2280;
defparam prom_inst_12.INIT_RAM_1B = 256'h8E57796AC8D96EDCB6DB36DF30342E39B99BF251E4D920971B660C96C466AE4B;
defparam prom_inst_12.INIT_RAM_1C = 256'hB26DCCCBCF7F9BF3DDFE2F6D6CD99D59FE76DB6EDB9EC9065B339B65E5331EAC;
defparam prom_inst_12.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF72BECDB6DB13;
defparam prom_inst_12.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_12.INIT_RAM_20 = 256'h07261C939265C00E132E01C265C03932E07265C0732B87D29AD9000040555004;
defparam prom_inst_12.INIT_RAM_21 = 256'hF3007327F97FC9FE4FF27FFFDFF64B37A436E01C9872439265C0E4C0E49C932E;
defparam prom_inst_12.INIT_RAM_22 = 256'hD8C48C80AC6320A588B2C4D89666DB11620AF98050C9116499B124CD9666C415;
defparam prom_inst_12.INIT_RAM_23 = 256'h6CC58C1050C6605E97E9D0BD193168241431820BD3A172CD04C641434120BC6E;
defparam prom_inst_12.INIT_RAM_24 = 256'hB349CC20BD3A17449A209A4C48293461920A68B8DCC58C2484C480AC613920B4;
defparam prom_inst_12.INIT_RAM_25 = 256'hC6831A61A046846311D1362124262082B149C9817A5FA742EA88B66125104482;
defparam prom_inst_12.INIT_RAM_26 = 256'h46B11A0111A0C4699868191A118C476846D0641A46831A011AC68386831AC680;
defparam prom_inst_12.INIT_RAM_27 = 256'h7C6C89B2C458B662D931620AF98073431B409106B11A0C4680C46991A0661A06;
defparam prom_inst_12.INIT_RAM_28 = 256'hD191A00EE6341C3405B428D83407311A011A02B226C93162488B6CCD882BE601;
defparam prom_inst_12.INIT_RAM_29 = 256'h40576850910680EE62340623405A502C680EE60D0234216858D007731A0C6C02;
defparam prom_inst_12.INIT_RAM_2A = 256'h7352941B223407311068311A10ACC8D0873191A0446C02D0B11A00EE32340CC3;
defparam prom_inst_12.INIT_RAM_2B = 256'hCD4646804680AC8D01DCE1A02970D01CD6851906811A00AC8D007711A0292340;
defparam prom_inst_12.INIT_RAM_2C = 256'h4246811A00AC8D007731A10A58D08735294191A041A02B20D01DCC6C02963601;
defparam prom_inst_12.INIT_RAM_2D = 256'h14911A03B88834056661A03B8DA142C41A0446802B323421DCE4680A5C8D01CD;
defparam prom_inst_12.INIT_RAM_2E = 256'h0852646843BA86940911A0C41A029620D01CC646C02B323601DD42588D0088D0;
defparam prom_inst_12.INIT_RAM_2F = 256'hF4596C4122C23839C896C4122D22BE6414B6FE84B2234188D0056C46C039888D;
defparam prom_inst_12.INIT_RAM_30 = 256'h6C35F6B73ECFB7DFD9F67D9F67D6C6C413211C1CE6362082CFB3EDF5FA9F67D9;
defparam prom_inst_12.INIT_RAM_31 = 256'h0E77E96C7D9F7F5FA8FB3EDF7F4865B04707395F4C900096C11C1CE5FA2562BE;
defparam prom_inst_12.INIT_RAM_32 = 256'h0470664D9225B8238332675BF8FB3EDF7F63ECFB7DFD646C11C1CE2C8263608E;
defparam prom_inst_12.INIT_RAM_33 = 256'h67D9F67DFD2096C110448C4B6088225FAFD16CFB3ECFB3EBF53ECFB3ECFA2CB7;
defparam prom_inst_12.INIT_RAM_34 = 256'hD9F5FA9F67D9F67D9F4C96C104707390932D8208E0E72652FE7D9F67D4FBFA9F;
defparam prom_inst_12.INIT_RAM_35 = 256'h4FBFAFD7EB04B60823839C48CCB608230207394FB3ECFB3ECFBFA2D9F67D9F67;
defparam prom_inst_12.INIT_RAM_36 = 256'h7D7EA7D325B0411C1839C84996C1046040E729F67D9F67D9F4B4BF9F67D9F67D;
defparam prom_inst_12.INIT_RAM_37 = 256'h2196C1047060E712712D8200C081CC013ECFB3ECFB3ECFBFA2D9F67D9F67D9F6;
defparam prom_inst_12.INIT_RAM_38 = 256'h3073890912D8200C081CC253ECFB3ECFB3ECFACADFCFB3ECFB3ECFA9F7F5FAFD;
defparam prom_inst_12.INIT_RAM_39 = 256'h001810398027D9F67D9F67D9F67DFD16CFB3ECFB3ECFB3ECFAFD4FA2CB608238;
defparam prom_inst_12.INIT_RAM_3A = 256'h7D9F67D9F67D652FE7D9F67D9F67D9F53EFEBF5FAC12D82088E0C1CE24665B00;
defparam prom_inst_12.INIT_RAM_3B = 256'hF67D9F67D9F67D9F67D7EA7D165B04111C1839C484896C00006040E60467D9F6;
defparam prom_inst_12.INIT_RAM_3C = 256'hAFD6096C104471060E712332D00000C0081CC013ECFB3ECFB3ECFB3ECFBFA2D9;
defparam prom_inst_12.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCFB3ECFB3ECFB3ECFA9F7F5F;
defparam prom_inst_12.INIT_RAM_3E = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000;
defparam prom_inst_12.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFF000000000000000000000000FFFFFFFFFFFFFFFF;

pROM prom_inst_13 (
    .DO({prom_inst_13_dout_w[30:0],prom_inst_13_dout[6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_13.READ_MODE = 1'b0;
defparam prom_inst_13.BIT_WIDTH = 1;
defparam prom_inst_13.RESET_MODE = "SYNC";
defparam prom_inst_13.INIT_RAM_00 = 256'hDB6DB6DB6D4591A9252083641231248054618836552AC883497FFFC2FFFF0087;
defparam prom_inst_13.INIT_RAM_01 = 256'hD064D90888A22228888A222333223222222248B22322222362C37284CEDB6DB6;
defparam prom_inst_13.INIT_RAM_02 = 256'h9556FBF0BB6DDF7DF5DB6EF700295463DED12E7D2ECB2A8888888888C88B79BC;
defparam prom_inst_13.INIT_RAM_03 = 256'h3022B22A60C9B383EB8C99121598C99121598C99121599B44C8D599B44C8D595;
defparam prom_inst_13.INIT_RAM_04 = 256'hDA2746AEC56632FA8ACF95958CC99999B344FB359B6DB6CDC624CB14D4D40DCB;
defparam prom_inst_13.INIT_RAM_05 = 256'hF49204558ADF6F8332222332D98D98D9876DC8C3FE4AD761AA045C936903CD6C;
defparam prom_inst_13.INIT_RAM_06 = 256'hFF2D57FCB55FF2E3FA56DF6FB8FE95CDA2646ACC5656CFF2CF15D3207FE9241F;
defparam prom_inst_13.INIT_RAM_07 = 256'h5865B7DBEFF3FFBAD7B5AF6EFFA326A0FBF7F56F4BEFB5FE5F7DAFF2D57FCB55;
defparam prom_inst_13.INIT_RAM_08 = 256'h956C7957577AE7DF58A5953B9ABABBB116EDE1807B116EDA1807BEFB71FFCBC4;
defparam prom_inst_13.INIT_RAM_09 = 256'h63BE98E149011384DB76FB7E748A9ADE6B53DBEDFED9FFFFFFF5E9903B298A98;
defparam prom_inst_13.INIT_RAM_0A = 256'hDE92E5CBDB7A5B7C32AD54F89CF6AB876D559E9912449E33718933CCC32C5225;
defparam prom_inst_13.INIT_RAM_0B = 256'h3DDFE32FDD8C88C8CCCCB6DB55DB6DEDB6DBDB6DBDB7A4B972F6DE92E5CB8F96;
defparam prom_inst_13.INIT_RAM_0C = 256'h83F49D35D2D23F9BEBD73B398F9CC7E73E2378E0C768D1078ABEAF73B9C7F9BF;
defparam prom_inst_13.INIT_RAM_0D = 256'h3B2E95FF3FBCF833BD35F73F69E09DE9FCDF5FB9D9EC7CF63F29F11BC7063398;
defparam prom_inst_13.INIT_RAM_0E = 256'hC5CFAE3437A493C0D0CB0E9A9D91131206428983A0209813BE25165165165165;
defparam prom_inst_13.INIT_RAM_0F = 256'hADDB68000000000090A42AAE55CB972AAAAAAB95572B0FDF303B75BD7B10965E;
defparam prom_inst_13.INIT_RAM_10 = 256'hDBB16FECBB6D8CC18CDFFB626EEDBBB771AB83666EEDBBB771AA0CD9B7FC8177;
defparam prom_inst_13.INIT_RAM_11 = 256'h08E236EC790B8FFEFEC9BA6D0B28C9117A27D1DFC04711B763C85C7C889B7DBE;
defparam prom_inst_13.INIT_RAM_12 = 256'h1DC238C338BEECB8F999BB2DB06C603DE1B2EC9BB198CF072D19222F44DA3BD8;
defparam prom_inst_13.INIT_RAM_13 = 256'hDFEAAFF4FF770F935DB765ADC2E9B5B76CCEF77C672122D6DDB33DC7CF7DB440;
defparam prom_inst_13.INIT_RAM_14 = 256'hAC755EA8FFAAEA23CF55F72EF4BA1C1B145DA577E71FF58E4B7FA9FAD7F53F52;
defparam prom_inst_13.INIT_RAM_15 = 256'hFE6DB74552929293C6A4689612D0B42D0BBD77342EB5D52492492CEB31276664;
defparam prom_inst_13.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF4B905294BCD2D55277A;
defparam prom_inst_13.INIT_RAM_17 = 256'h0000FFFFFFFFFFFFFFFF000000000000FFFFF7C0FFFFFC7C3D3133FE38FFFE38;
defparam prom_inst_13.INIT_RAM_18 = 256'h00000000000000000000FFFFFFFFFFFF000003FF000103E7FFFFFC0F00000000;
defparam prom_inst_13.INIT_RAM_19 = 256'hFFFFFAABFFABFEAFAAAAAAAAAAEAFEBAAAAAAAAAAABAFABBAAAAAAAAEEAAAAAA;
defparam prom_inst_13.INIT_RAM_1A = 256'h2A82882A80AFBDE083BB33F92FD65820576F76C10362D9040ABADA9202272BEE;
defparam prom_inst_13.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000AAAAAA0002AA02A82A08288A208A0;
defparam prom_inst_13.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_13.INIT_RAM_20 = 256'h441504551510555F55554000154015014141044444140005110011004040417F;
defparam prom_inst_13.INIT_RAM_21 = 256'h5041441104505540445541415045144F55555000154015415041444144501501;
defparam prom_inst_13.INIT_RAM_22 = 256'h55555000155005415051441114505550445011004540000F5555500015500541;
defparam prom_inst_13.INIT_RAM_23 = 256'h110541404545150F55555000155005405051451110415554114004551015410F;
defparam prom_inst_13.INIT_RAM_24 = 256'h5050411111454005041551151010150F55555000155005405050451111415015;
defparam prom_inst_13.INIT_RAM_25 = 256'h55555000155005405050411111050001445014554545405F5555500015500540;
defparam prom_inst_13.INIT_RAM_26 = 256'h105411545441557E5555000055005405050411111050001444004401010105FE;
defparam prom_inst_13.INIT_RAM_27 = 256'h4105104411415501115505054114513E55554000550055054105110511405405;
defparam prom_inst_13.INIT_RAM_28 = 256'h55554000554015054145104451415541114044011500003F5555400055401505;
defparam prom_inst_13.INIT_RAM_29 = 256'h441505011514543F55554000554015014145144441055550450011544055043F;
defparam prom_inst_13.INIT_RAM_2A = 256'h4141044445150014105544544040543F55554000554015014141144445054054;
defparam prom_inst_13.INIT_RAM_2B = 256'h55554000554015014141044444140005114051551515017F5555400055401501;
defparam prom_inst_13.INIT_RAM_2C = 256'h4514155411141440000000055555540005540550541051144114055011055055;
defparam prom_inst_13.INIT_RAM_2D = 256'h0554015014145144441055550450051500000001555554000554015054145104;
defparam prom_inst_13.INIT_RAM_2E = 256'h0000000155555400055401501414514444105415044141100000000155555400;
defparam prom_inst_13.INIT_RAM_2F = 256'h4441400051150515000000015555540005540150141411444451500145455441;
defparam prom_inst_13.INIT_RAM_30 = 256'h0554015014141044444140005110011000000001555554000554015014141044;
defparam prom_inst_13.INIT_RAM_31 = 256'h0000000155555400055401501404104414410050105050410000000155555400;
defparam prom_inst_13.INIT_RAM_32 = 256'h1450555044505100000000155555500015501541504144510450154044154155;
defparam prom_inst_13.INIT_RAM_33 = 256'h1550054050514511104155541140145500000005555550001550054150514411;
defparam prom_inst_13.INIT_RAM_34 = 256'h0000000555555000155005405051451110415054110504400000000555555000;
defparam prom_inst_13.INIT_RAM_35 = 256'h1105000144541455000000055555500015500540505045111145400515155104;
defparam prom_inst_13.INIT_RAM_36 = 256'h1550054050504111110500014440044000000005555550001550054050504111;
defparam prom_inst_13.INIT_RAM_37 = 256'h0000000555555000155005405010411051040140414141050000000555555000;
defparam prom_inst_13.INIT_RAM_38 = 256'h5555400000000000155555555555400000000000555555555555000000000000;
defparam prom_inst_13.INIT_RAM_39 = 256'h0000000001555555555554000000000005555555555550000000000005555555;
defparam prom_inst_13.INIT_RAM_3A = 256'h0015555555555540000000000055555555555500000000000055555555555400;
defparam prom_inst_13.INIT_RAM_3B = 256'h5555555400000000000555555555555000000000000555555555554000000000;
defparam prom_inst_13.INIT_RAM_3C = 256'h4000000000005555555555550000000000005555555555540000000000015555;
defparam prom_inst_13.INIT_RAM_3D = 256'h0000055555555555500000000000055555555555400000000000155555555555;
defparam prom_inst_13.INIT_RAM_3E = 256'h5555555555000000000000555555555554000000000001555555555554000000;
defparam prom_inst_13.INIT_RAM_3F = 256'h5550000000000005555555555540000000000015555555555540000000000055;

pROM prom_inst_14 (
    .DO({prom_inst_14_dout_w[30:0],prom_inst_14_dout[7]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_14.READ_MODE = 1'b0;
defparam prom_inst_14.BIT_WIDTH = 1;
defparam prom_inst_14.RESET_MODE = "SYNC";
defparam prom_inst_14.INIT_RAM_00 = 256'hFFFFFFFFFFC000000000000000000000FCC5457FFFFFBD000AF9FFFFFFFFFF83;
defparam prom_inst_14.INIT_RAM_01 = 256'h531AA341A270580CA5722E12D2C9570011B2555511001B000000000000000000;
defparam prom_inst_14.INIT_RAM_02 = 256'hFFFFFFFFFFFEBBB6D82B220398A57EA0D55042D951B4AFF104470E1C3A62AAAB;
defparam prom_inst_14.INIT_RAM_03 = 256'h14292D4A0945204A294945254AAD2AA2400092A5001054000000140050045550;
defparam prom_inst_14.INIT_RAM_04 = 256'h6AD66D6B76D6A3A120154B2080B9161A801548C4310C405251414312902B1295;
defparam prom_inst_14.INIT_RAM_05 = 256'h4B58ACACACACA564A498D4D43512521B50DA8C99144450B312954AA4AC4A57B3;
defparam prom_inst_14.INIT_RAM_06 = 256'hFFFFFFFFFFFFFFFEAA552957A952A7A96A551504862524A8949894A8C4918989;
defparam prom_inst_14.INIT_RAM_07 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5251B946EA4A36A5;
defparam prom_inst_14.INIT_RAM_0A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_0B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_0C = 256'h8888888C8980512A492544D39D269CE9552882A97A73A608915498A518249552;
defparam prom_inst_14.INIT_RAM_0D = 256'h154A4EF492769249312200635091300483B00724888C244446122232CCC88C88;
defparam prom_inst_14.INIT_RAM_0E = 256'h32484A24C90824C92554552932C924964924921212D5455293925544A4AA4955;
defparam prom_inst_14.INIT_RAM_0F = 256'h534E88B41A890A04C2B17F85055956618C60542BE0150020A18C40552898A933;
defparam prom_inst_14.INIT_RAM_10 = 256'h4A49E49E59254CC91C2528ADE4896AA5464D2751CD19824902400055035031C0;
defparam prom_inst_14.INIT_RAM_11 = 256'hDC10001010002018000804104C0810008104035123AA4C960B0592532A49E092;
defparam prom_inst_14.INIT_RAM_12 = 256'hE12196C21513A068DCB2084011E3333BB2ECBB22242108420421196484223C4D;
defparam prom_inst_14.INIT_RAM_13 = 256'h12A0ABD11168A2DA8AFA0029F40053F400A7E8014F68029E68053C340A7800C1;
defparam prom_inst_14.INIT_RAM_14 = 256'h16B00084A2095F4445A28B03FF18F4445A311F4445A28589FFFFFFFE3088022D;
defparam prom_inst_14.INIT_RAM_15 = 256'h3E6C03C989B2492492636692644E5CA0924929A235528A8935255288888B1D11;
defparam prom_inst_14.INIT_RAM_16 = 256'hFFFFFFF9AAA35300000004010184C4093102408124671332492663189CE4A925;
defparam prom_inst_14.INIT_RAM_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_18 = 256'hAAAAAA8000000002AAAAAA00000AAAA0002AA002A802A0A82820000008800000;
defparam prom_inst_14.INIT_RAM_19 = 256'h0000000002AAAAAAAAAAAAAAAAAAAAAAAAAAAAAA0000000000000000002AAAAA;
defparam prom_inst_14.INIT_RAM_1A = 256'h02008516C0000AC9D00C176A62244040208E354AABE015000200208000002080;
defparam prom_inst_14.INIT_RAM_1B = 256'h0443313F80512E489249924F1090041110C9F2D125A960B209404CB26407FC01;
defparam prom_inst_14.INIT_RAM_1C = 256'hA91AA2A52F6FECFDE6F93DE5264CBFF1FEF24926491C490C4962C940E9620FF8;
defparam prom_inst_14.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF68AA6C924911;
defparam prom_inst_14.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_14.INIT_RAM_20 = 256'h252A94B294ACC10A15660942ACC429566252ACC4C1398E00CA09000055015555;
defparam prom_inst_14.INIT_RAM_21 = 256'h5108236C7B23D91EC8F6C7FA48F64B3602226214AA52C294ACC4A550A594A566;
defparam prom_inst_14.INIT_RAM_22 = 256'hDCACD9820E56620598A644D096629911421AA890D04B134C89A164CD16628435;
defparam prom_inst_14.INIT_RAM_23 = 256'h66EDD8010AECE10A89A9504D09BB700C42BB002152A092E601ACC42980621452;
defparam prom_inst_14.INIT_RAM_24 = 256'h19CB0802152A090CDC20165A5881B84096206828A584DA2DC5858206D1616214;
defparam prom_inst_14.INIT_RAM_25 = 256'h4109046042410C6311D01731672C2008398B4B842A26A5412281B3396E100588;
defparam prom_inst_14.INIT_RAM_26 = 256'h411905099042641198109904318C436846D06404410B040904C10B010B044142;
defparam prom_inst_14.INIT_RAM_27 = 256'h54AD98A644D0B2228933421AA884A3071B41910131042C4102C4131042C4042C;
defparam prom_inst_14.INIT_RAM_28 = 256'h50904098F2084C084CB42858084C79040904263222991142C98A2C4D086AA213;
defparam prom_inst_14.INIT_RAM_29 = 256'h84C768519101098F2208122084CA50241098760216086328C8210C3904241426;
defparam prom_inst_14.INIT_RAM_2A = 256'hC3D2941962084C791010B104218D88210C7B1042E41426519904098772085CC0;
defparam prom_inst_14.INIT_RAM_2B = 256'h0F42410241098C82131EE04263702131F6851B010B0421858210C3B042616084;
defparam prom_inst_14.INIT_RAM_2C = 256'h46410904098C8204C7B04318D8218C7D2941B042C04261602130E41426120A13;
defparam prom_inst_14.INIT_RAM_2D = 256'h309904263CCC084C66604263DDA142C404244108612208430EC410985882130F;
defparam prom_inst_14.INIT_RAM_2E = 256'h18C26410C63E8E94091042C4042636202131EC414261620A130F46C88204C821;
defparam prom_inst_14.INIT_RAM_2F = 256'hD4D9100202C4106A819100206D26AA249CD6EA8DB2208488204C26410261CC82;
defparam prom_inst_14.INIT_RAM_30 = 256'h2CBD57BB1AC6B35B58D6358D635241002362083542080106C6B1ACD56A8D6358;
defparam prom_inst_14.INIT_RAM_31 = 256'h1AB5A92C358D6D56A86B1ACD6D482440830D504D4D808091020835656A2D66AA;
defparam prom_inst_14.INIT_RAM_32 = 256'h0820A805806460410540654BA86B1ACD6D61AC6B35B564102083546404608104;
defparam prom_inst_14.INIT_RAM_33 = 256'h6358D635B5699102008018C881004256AB536C6B1AC6B1AAD51AC6B1AC6A6C8C;
defparam prom_inst_14.INIT_RAM_34 = 256'h58D56A8D6358D6358D4591020820D5000122041041AA02D2EA358D63546B6A8D;
defparam prom_inst_14.INIT_RAM_35 = 256'h46B6AB55A90C88104106A801848A1861870D5946B1AC6B1AC6B6A6D8D6358D63;
defparam prom_inst_14.INIT_RAM_36 = 256'h355AA35164408208306A800091430C30E1AA08D6358D6358D5B4BA8D6358D635;
defparam prom_inst_14.INIT_RAM_37 = 256'h6191020820C1AA006322861861C356251AC6B1AC6B1AC6B6A6D8D6358D6358D6;
defparam prom_inst_14.INIT_RAM_38 = 256'h60D50000322861861C356011AC6B1AC6B1AC6ACA5D46B1AC6B1AC6A8D6D56AB5;
defparam prom_inst_14.INIT_RAM_39 = 256'h310C386AC4A358D6358D6358D635B512C6B1AC6B1AC6B1AC6AB546A6C8810410;
defparam prom_inst_14.INIT_RAM_3A = 256'h358D6358D6352D2EA358D6358D6358D51ADAAD56AC122041004183540046450C;
defparam prom_inst_14.INIT_RAM_3B = 256'hD6358D6358D6358D6355AA351244082008306A8000091430C430E1AB0CE358D6;
defparam prom_inst_14.INIT_RAM_3C = 256'hAB5219102080200C1AA00612286188621C356251AC6B1AC6B1AC6B1AC6B6A6D8;
defparam prom_inst_14.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFC6B1AC6B1AC6B1AC6A8D6D56;
defparam prom_inst_14.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFF000000000000000000000000000000000000000000000000;
defparam prom_inst_14.INIT_RAM_3F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000;

pROM prom_inst_15 (
    .DO({prom_inst_15_dout_w[30:0],prom_inst_15_dout[7]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD(ad[13:0])
);

defparam prom_inst_15.READ_MODE = 1'b0;
defparam prom_inst_15.BIT_WIDTH = 1;
defparam prom_inst_15.RESET_MODE = "SYNC";
defparam prom_inst_15.INIT_RAM_00 = 256'h4924924924614A249091800C006012025C049C0055000143217FFFC2FFFF3447;
defparam prom_inst_15.INIT_RAM_01 = 256'h5152010888A22228888A22223223222222220CA232222223626122028A492492;
defparam prom_inst_15.INIT_RAM_02 = 256'h5506AAAAA5A44B55552D225280255661CED16C35A6DB88088888888888893098;
defparam prom_inst_15.INIT_RAM_03 = 256'h6822A92D50A551454B5A54285555A54285555A54285559B00A05559B00A05555;
defparam prom_inst_15.INIT_RAM_04 = 256'hD80402A8A5556AA34AAE15555AA89911BB00F0000000001000122A947A7A2D23;
defparam prom_inst_15.INIT_RAM_05 = 256'h46DBC4554E4F2783332232324B44B44B4524A580FD2AD751AB345A4924A30D6C;
defparam prom_inst_15.INIT_RAM_06 = 256'hFEA553FA954FEA417D164F27905F45CD80502AAA5556AFEAAE9768917C8DB79E;
defparam prom_inst_15.INIT_RAM_07 = 256'h492193C9FBF9EABEF6B5AFBAAAA423D12A54A54D49A695FD4D34AFEA553FA954;
defparam prom_inst_15.INIT_RAM_08 = 256'h416AF554547AE5D7500715A182A2A391126CA304B91126CA104B9E7920BF43C4;
defparam prom_inst_15.INIT_RAM_09 = 256'h833410406D3E1184D932793C3C88129A7A03C9E4FA48FEFCAAA5B448BB2D8815;
defparam prom_inst_15.INIT_RAM_0A = 256'h4E964C99C93A493A6BAF40E8357FA913FF441D44390E546123554BC9890C0255;
defparam prom_inst_15.INIT_RAM_0B = 256'hDE6F56AFDDC88888CCCC924955C924E49249C9249C93A59326724E964C990792;
defparam prom_inst_15.INIT_RAM_0C = 256'h0574DD1993925EEABBF71F214790A3E52D0479A18A91220A82BEAFD3E9E4FECF;
defparam prom_inst_15.INIT_RAM_0D = 256'h3C885CFD2AFCA82A153CFD29F92050A9FF55DEB8D92A3C951F296823CD0C5601;
defparam prom_inst_15.INIT_RAM_0E = 256'h34CF2D7A022AABA0682AA69A0D12A931452398221051552AE812924904124904;
defparam prom_inst_15.INIT_RAM_0F = 256'hB1382C000000000090A42AAB556AD5AAAAAAAAD555AA83062A29349D20D0D748;
defparam prom_inst_15.INIT_RAM_10 = 256'h499127AC3A648440864FA927666C9B9370E38123666C9B9370E2064893EA8077;
defparam prom_inst_15.INIT_RAM_11 = 256'h08A2225E65891EF7DE599A24031888012622B08AC0451112F32C48F888D93C9E;
defparam prom_inst_15.INIT_RAM_12 = 256'h11026011A436E5906021B96490B83030B093E599B0B05D920F110024C4561158;
defparam prom_inst_15.INIT_RAM_13 = 256'h9F7AA7BE7BD32E105E372CF142FA1CF26C6E453003212673C9B1BDF70F300022;
defparam prom_inst_15.INIT_RAM_14 = 256'hAC7552A97FAAEA211815750FF43F302F0849A5D9B214D88A093DF5DF17BEBBEA;
defparam prom_inst_15.INIT_RAM_15 = 256'hFE60000553838383C7A4A902024090240B2D65102CB5972090482CAB21041E65;
defparam prom_inst_15.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF53984210BCC2155077A;
defparam prom_inst_15.INIT_RAM_17 = 256'h00000000000000000000FFFF0000000000000BDF00000067843DC00F07FFFFC0;
defparam prom_inst_15.INIT_RAM_18 = 256'h00000000000000000000FFFFFFFFFFFF000003FF000103E7FFFFFC0F00000000;
defparam prom_inst_15.INIT_RAM_19 = 256'hFFFFFAABFFFEAAAFAFAEAAAABFBEAAAAAAAAAAAAAAAAFEEBAAAAAAAAEFEAAAAA;
defparam prom_inst_15.INIT_RAM_1A = 256'hA208A02A828D1EE104E089D8B59A684104F7A242089B8B08222A48DA7C2321AE;
defparam prom_inst_15.INIT_RAM_1B = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFF80000000000000AAAAAA0002AA02A82A08288;
defparam prom_inst_15.INIT_RAM_1C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_1F = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam prom_inst_15.INIT_RAM_20 = 256'h5015014415045515000015555540005540150141410444441400051100110040;
defparam prom_inst_15.INIT_RAM_21 = 256'h5015415041441104505540445541415000000555554000155015414041445144;
defparam prom_inst_15.INIT_RAM_22 = 256'h0000055555500015500541505144111450555044501100450000055555500015;
defparam prom_inst_15.INIT_RAM_23 = 256'h4150151105414045000005555550001550054050514511104155541140045510;
defparam prom_inst_15.INIT_RAM_24 = 256'h5005405050411111454005041551151000000555555000155005405050451111;
defparam prom_inst_15.INIT_RAM_25 = 256'h0000055555500015500540505041111105000144501455450000055555500015;
defparam prom_inst_15.INIT_RAM_26 = 256'h4054051054115454000055555500015500540505041111105000144400440101;
defparam prom_inst_15.INIT_RAM_27 = 256'h4055054105104411415501115505054100001555550000554055050105114511;
defparam prom_inst_15.INIT_RAM_28 = 256'h0000155555400055401505414510445141554111404401150000155555400055;
defparam prom_inst_15.INIT_RAM_29 = 256'h0540544415050115000015555540005540150141451444410555504500115440;
defparam prom_inst_15.INIT_RAM_2A = 256'h4015014141044445150014105544544000001555554000554015014141144445;
defparam prom_inst_15.INIT_RAM_2B = 256'h0000155555400055401501414104444414000511405155150000155555400055;
defparam prom_inst_15.INIT_RAM_2C = 256'h1451044514155411000000000000015555540005540550541051144114055011;
defparam prom_inst_15.INIT_RAM_2D = 256'h5554000554015014145144441055550400000000000001555554000554015054;
defparam prom_inst_15.INIT_RAM_2E = 256'h0000000000000155555400055401501414514444105415040000000000000155;
defparam prom_inst_15.INIT_RAM_2F = 256'h1410444441400051000000000000015555540005540150141410444451500145;
defparam prom_inst_15.INIT_RAM_30 = 256'h5554000554015014141044444140005100000000000001555554000554015014;
defparam prom_inst_15.INIT_RAM_31 = 256'h0000000000000155555400055401501404104414410050100000000000000155;
defparam prom_inst_15.INIT_RAM_32 = 256'h5144111450555044000000000000055555500015501541504144510450154044;
defparam prom_inst_15.INIT_RAM_33 = 256'h5550001550054050514511104155541100000000000005555550001550054150;
defparam prom_inst_15.INIT_RAM_34 = 256'h0000000000000555555000155005405051451110415054110000000000000555;
defparam prom_inst_15.INIT_RAM_35 = 256'h5041111105000144000000000000055555500015500540505041111145400515;
defparam prom_inst_15.INIT_RAM_36 = 256'h5550001550054050504111110500014400000000000005555550001550054050;
defparam prom_inst_15.INIT_RAM_37 = 256'h0000000000000555555000155005405010411051040140410000000000000555;
defparam prom_inst_15.INIT_RAM_38 = 256'h0000000000000000155555555555555555555555000000000000000000000000;
defparam prom_inst_15.INIT_RAM_39 = 256'h5555555554000000000000000000000005555555555555555555555550000000;
defparam prom_inst_15.INIT_RAM_3A = 256'h0015555555555555555555555500000000000000000000000055555555555555;
defparam prom_inst_15.INIT_RAM_3B = 256'h0000000000000000000555555555555555555555555000000000000000000000;
defparam prom_inst_15.INIT_RAM_3C = 256'h5555555555550000000000000000000000005555555555555555555555540000;
defparam prom_inst_15.INIT_RAM_3D = 256'h0000055555555555555555555555500000000000000000000000155555555555;
defparam prom_inst_15.INIT_RAM_3E = 256'h0000000000000000000000555555555555555555555554000000000000000000;
defparam prom_inst_15.INIT_RAM_3F = 256'h5555555555555550000000000000000000000015555555555555555555555500;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[14]),
  .CLK(clk),
  .CE(ce)
);
MUX2 mux_inst_0 (
  .O(dout[0]),
  .I0(prom_inst_0_dout[0]),
  .I1(prom_inst_1_dout[0]),
  .S0(dff_q_0)
);
MUX2 mux_inst_1 (
  .O(dout[1]),
  .I0(prom_inst_2_dout[1]),
  .I1(prom_inst_3_dout[1]),
  .S0(dff_q_0)
);
MUX2 mux_inst_2 (
  .O(dout[2]),
  .I0(prom_inst_4_dout[2]),
  .I1(prom_inst_5_dout[2]),
  .S0(dff_q_0)
);
MUX2 mux_inst_3 (
  .O(dout[3]),
  .I0(prom_inst_6_dout[3]),
  .I1(prom_inst_7_dout[3]),
  .S0(dff_q_0)
);
MUX2 mux_inst_4 (
  .O(dout[4]),
  .I0(prom_inst_8_dout[4]),
  .I1(prom_inst_9_dout[4]),
  .S0(dff_q_0)
);
MUX2 mux_inst_5 (
  .O(dout[5]),
  .I0(prom_inst_10_dout[5]),
  .I1(prom_inst_11_dout[5]),
  .S0(dff_q_0)
);
MUX2 mux_inst_6 (
  .O(dout[6]),
  .I0(prom_inst_12_dout[6]),
  .I1(prom_inst_13_dout[6]),
  .S0(dff_q_0)
);
MUX2 mux_inst_7 (
  .O(dout[7]),
  .I0(prom_inst_14_dout[7]),
  .I1(prom_inst_15_dout[7]),
  .S0(dff_q_0)
);
endmodule //rom_gs105b
