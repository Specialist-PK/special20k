//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.11 (64-bit)
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Tue Apr  8 22:07:07 2025

module t20k_rom (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [12:0] ad;

wire [29:0] prom_inst_0_dout_w;
wire [29:0] prom_inst_1_dout_w;
wire [29:0] prom_inst_2_dout_w;
wire [29:0] prom_inst_3_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[29:0],dout[1:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 2;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'hE552E0B2CBC8D6F83577E2D9F6E2A8C82655557A2935555C7A07A41500FEAF4F;
defparam prom_inst_0.INIT_RAM_01 = 256'h9A27A9E6589E2499EA78B21F2041252C2CBA09959B4EFAD55095DDCDD9C88A74;
defparam prom_inst_0.INIT_RAM_02 = 256'hA77EED9518E7B6CBC8104017E96657E966597F96A1727C957E966497F9EA177B;
defparam prom_inst_0.INIT_RAM_03 = 256'hD7CB2696F9AADA15E6E2E9EECA9BAB685AF2B795FE551D89BD4595495546977E;
defparam prom_inst_0.INIT_RAM_04 = 256'hE5169BBB687B62F97E67EA5D1C958B4BFDBB1860A5EF65EA66EEDA1E6A4EEE3E;
defparam prom_inst_0.INIT_RAM_05 = 256'hBE7EF246FB2E991E8A157AE1B5BD0FC955564FA55CBF287B2FC8FBD5647D5D96;
defparam prom_inst_0.INIT_RAM_06 = 256'hB6C940004A225209FC13A3CBE5F94789561563763EBDF8A3476ACB22CBE172AC;
defparam prom_inst_0.INIT_RAM_07 = 256'hBF780157A41F9B07FA9BE2D54FF957EE96FBBA6CFEFAA7AEDB6D77ED8A2DBF9D;
defparam prom_inst_0.INIT_RAM_08 = 256'h0020021DB7EF8EA09BD7ED4117D04D0F342E4637E9D20BE42CDFD2FD2FD2FBF4;
defparam prom_inst_0.INIT_RAM_09 = 256'h00CEE4E40044E4E70089F9DE0088387600F0817900600D91316F83000CFA0C1A;
defparam prom_inst_0.INIT_RAM_0A = 256'h0024000000C0000000C0019002A02002002A19283C24098C2BBA002A00000000;
defparam prom_inst_0.INIT_RAM_0B = 256'h00960260033020020000000009D625960027258325632BAA25A7309620002576;
defparam prom_inst_0.INIT_RAM_0C = 256'h25561755155D340018092555200215D537060083308325562406259617582376;
defparam prom_inst_0.INIT_RAM_0D = 256'hC00000182AAA0600200230A70025162525550295255500032586189619560096;
defparam prom_inst_0.INIT_RAM_0E = 256'h255615D5155D15571C0D1575157516250007035C32A31EAA1EAA258317562556;
defparam prom_inst_0.INIT_RAM_0F = 256'hFFFF15D51D5525D6355525961555258025961595009520072406009615D71557;
defparam prom_inst_0.INIT_RAM_10 = 256'hA9EE288E22B86259AE217D565E4B37EB7607D2CB0477D30638E79E3EF38FFFCB;
defparam prom_inst_0.INIT_RAM_11 = 256'h76441F9107644A5752E717E7E415FEFE50547E50BA38BB6E2A92E698AA188AE4;
defparam prom_inst_0.INIT_RAM_12 = 256'h9F6FB6F41F9765FBD9AF4B757114799579076EBED5B9AF779657655465117B90;
defparam prom_inst_0.INIT_RAM_13 = 256'h6971979071C5E5E6F4A9E6F7BECB9C75975F9AD8FA8B5F90556BFAAD2D145907;
defparam prom_inst_0.INIT_RAM_14 = 256'h72526F5971AC1CA5D41FA5E41EA5C7D88D1E85FBCBEBF4BF4B5BFEADE6B5C6AF;
defparam prom_inst_0.INIT_RAM_15 = 256'hAFC8DC6C6C7C4C55C6B9E79AFC6AEC6A716EC6B9EA2D4B9B6B1E71C65D7E4155;
defparam prom_inst_0.INIT_RAM_16 = 256'h656D9726CF8A2C55F361287A127C97A0CF61DF6C8DDBE6C8BD472712EAF1317E;
defparam prom_inst_0.INIT_RAM_17 = 256'hF7A65ED0F6171E9C1CB6F07A7D957E77ACE6E9BCB69435EB97A557F1F9147E57;
defparam prom_inst_0.INIT_RAM_18 = 256'h14559656512FC35F65965965814EA3FC368BC352F0D7D965604A659656DF7755;
defparam prom_inst_0.INIT_RAM_19 = 256'hF87647E47647CAC47F652B43658686E389D0BDA2055DF18D0C1E138D76050597;
defparam prom_inst_0.INIT_RAM_1A = 256'h520E1F499E2000000079BDC51715227A2E89B92A889DFF555D58868172DBF876;
defparam prom_inst_0.INIT_RAM_1B = 256'h8BA26E9AA62519F7FF67D5753D3F55625AA9F659607DF5574E1287A12D236749;
defparam prom_inst_0.INIT_RAM_1C = 256'hFB8B8BAABB2A5561652CEF4E86FF658B43659620584A7E10BA7975498749E61D;
defparam prom_inst_0.INIT_RAM_1D = 256'hB6EABAA53642C9656529798890E54BA6AE787E1FFD5878695639BBB685B93BB9;
defparam prom_inst_0.INIT_RAM_1E = 256'h8000011157160E2F0CB1B4A179F18696165A29572076727F2EBE7FBF88890552;
defparam prom_inst_0.INIT_RAM_1F = 256'h04C7050121041441C618500024FC6079F9136109A6F84D849819A089A0C49854;
defparam prom_inst_0.INIT_RAM_20 = 256'h7B6ECFF0BE388EE3FC2A2BA97BA541069065645A05106519CA926421F2C51049;
defparam prom_inst_0.INIT_RAM_21 = 256'hA54AE6D16C5BA4B06518A1481E14812189934EE351B9A42CA2B84998BF34245E;
defparam prom_inst_0.INIT_RAM_22 = 256'h439455CD6AAA6A188296D6B268A8461610690410E90DA4394E70D1B5ADA2BB43;
defparam prom_inst_0.INIT_RAM_23 = 256'h369AC5151445245451FE3EEEE45690534105EAB7BADE6B56A9185A5D85E56A9B;
defparam prom_inst_0.INIT_RAM_24 = 256'hAA2E2058AD2AB62A81D6279E288AA7AF5996E5F148521496A5717F18AA29BA62;
defparam prom_inst_0.INIT_RAM_25 = 256'h4628F85163624070CC90E4FA21A47C7118E264941A5E36655FA6E99A6A98A220;
defparam prom_inst_0.INIT_RAM_26 = 256'hAF5B66E4991BD297A712A56C931EF9841E5BEE2797939F9B95C410508315402E;
defparam prom_inst_0.INIT_RAM_27 = 256'hE2A85D4D57E4A1ABB9E797E4A1E79E7A2E7DAE9B560412BDEDAB9E79E5F66F58;
defparam prom_inst_0.INIT_RAM_28 = 256'h5D286E2B9971C4E79EE78B9A72D4B2E571C4E7F9FE48A75D72D5B2E5493D5F24;
defparam prom_inst_0.INIT_RAM_29 = 256'h6BCAF01FFF40004C30D5151519CD0457CF7EFDCBDBEBF9CBDBEBF9BBB9F22604;
defparam prom_inst_0.INIT_RAM_2A = 256'h2DA489EE549F24B92A7A9AD1E78E1A7FCF97CF19593F294949FE12D05C356EEE;
defparam prom_inst_0.INIT_RAM_2B = 256'h78BA8B44704F50D17BE11B4AB4BA179E7C8B7B934AA779DA924BA5EA23474F6F;
defparam prom_inst_0.INIT_RAM_2C = 256'h14A6A991611697481AA9A6A6E89616186ACDDDD89616146A549ADA16145A3044;
defparam prom_inst_0.INIT_RAM_2D = 256'hE60E10E1527EEE96262A49962CBCBCBDA525D9617624659B896E9BF66EA2EEE5;
defparam prom_inst_0.INIT_RAM_2E = 256'hE45B907B1595E9A3DC9EC918566E2DD969EEA765869CB595C5559BD882F21C7E;
defparam prom_inst_0.INIT_RAM_2F = 256'hFB9772F88ED2F88AFAABEAAFBBE4537BE9F547FF64D767957EF22FAE4ED6F8A6;
defparam prom_inst_0.INIT_RAM_30 = 256'h6D979AE1D4615B81465866C6E850A856799454B94A4424B9118B37BE5F4E6E05;
defparam prom_inst_0.INIT_RAM_31 = 256'h000000000000000000000000000000000000F51A56E0539A56E84EA1464B911E;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[29:0],dout[3:2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 2;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'h8EA1E27847F7C7C72AB761E2BC103FF8639560B600A555503A03480505303F00;
defparam prom_inst_1.INIT_RAM_01 = 256'hCAF1ACAB3AC6B2BC2B18FE03C2030F231F3911F8E78C7AE0031D439438EA4444;
defparam prom_inst_1.INIT_RAM_02 = 256'hB3F0BC952C2BFACCF080C00CE4C7CCE4E3F4C44A3CC1103CCE407C4C440FCC1B;
defparam prom_inst_1.INIT_RAM_03 = 256'hC4D3E2123401C87104F1C8CFC8B28721C2760F540F603C0D100D5A01600113F0;
defparam prom_inst_1.INIT_RAM_04 = 256'h8C3523C721FC23F9B03B03103D20D745561BFC811E5F210044F1C87D8ABBF48D;
defparam prom_inst_1.INIT_RAM_05 = 256'h86BE7663F3020C338C30F8C30C7802FA55801FA58F2BE3FFC0F9B78603786FA0;
defparam prom_inst_1.INIT_RAM_06 = 256'h724D40008C83218C2002C0CBC8030F4E00B5482C8E3C13C80C2BD3C1F80202BF;
defparam prom_inst_1.INIT_RAM_07 = 256'hF1FC02004DBC0E6FC3456B5501FA0B2019C3C0B330C078C6C722F0685A3CB76C;
defparam prom_inst_1.INIT_RAM_08 = 256'h020800EC88FF1EB8BC7B22DB7FC510601E3F9C5C0EB2D4F941747B47BC7BC11E;
defparam prom_inst_1.INIT_RAM_09 = 256'h00FA550000CA550200AB9D9200F5F01900FC26CC00E88AAC330703E0033E0C06;
defparam prom_inst_1.INIT_RAM_0A = 256'h02403C0000C027C005D405D4240606A4004531E9024A1DDD2BBA002A11550000;
defparam prom_inst_1.INIT_RAM_0B = 256'h110324060330062427CF3C3C30C330C32A4330C93033032430433243355D3243;
defparam prom_inst_1.INIT_RAM_0C = 256'h300300600058300001903000355700C0300300C330C33AAB300330C303093143;
defparam prom_inst_1.INIT_RAM_0D = 256'hC0000009300300603AAB32C315600260254016803000155730C301C3310300C3;
defparam prom_inst_1.INIT_RAM_0E = 256'h340700C000582AA901900241024002600003175D30C30EA90C0030C3030305D4;
defparam prom_inst_1.INIT_RAM_0F = 256'hFFFF00C00D55304335543043258030C030C305D409803557300300C309C30003;
defparam prom_inst_1.INIT_RAM_10 = 256'h8EA79AFA7EAFEFDBFE7CF3EFFC24AF8F3083C82C0B8A200ACF3CF3CA00E04124;
defparam prom_inst_1.INIT_RAM_11 = 256'hF6AFFDABFFEAECC8D7D34BAB8BF81EFBBFE6C378FF48BE23C9E678AF6FAAF638;
defparam prom_inst_1.INIT_RAM_12 = 256'h87ADB4080C0701F2F230A49C22BAC6BB38238DF4989AC6A0FFB6BF8AFFAB6E6F;
defparam prom_inst_1.INIT_RAM_13 = 256'h2FF0FFC5F0C28E8B1ECE8B1FF0C6BC30FF0F2A7A3CA98C23B568F2A792BAEB23;
defparam prom_inst_1.INIT_RAM_14 = 256'hBE8DDC1FFC83FFBFE3FCBFD3FEBFC33B172EBBCAF2E11EF1ECBA02A68AF0C2A7;
defparam prom_inst_1.INIT_RAM_15 = 256'h808970F0E0E0F0F00DEFBEF900E27C28C3B30DEFF22606B0FF0AF0C3FC308ED5;
defparam prom_inst_1.INIT_RAM_16 = 256'hA03E2E8F3B3F3C166C3BBEFFBB6BAE8BB03BD76B97D2EF8AC7DA0C33F803C3F2;
defparam prom_inst_1.INIT_RAM_17 = 256'hCE4F7FF07ABF4B13F57AAFECEE956043C34BF9DC3AFE5CF38788003CE3EDF656;
defparam prom_inst_1.INIT_RAM_18 = 256'h07B8EFFFFDD025CCFFFE4EFFFF72EE025CF025CD09733FFF7FFAB8EFF7B02C00;
defparam prom_inst_1.INIT_RAM_19 = 256'hD0B4CF0CF0CCC2C3CCFFC065FBEFFAFD8ECF9DB1FE220E17F3378E977302FCFF;
defparam prom_inst_1.INIT_RAM_1A = 256'hF4B3BDCBF6B0000000C8C7C17706119747D8F76BD8E3036ABBEBEF80B2CAC9F6;
defparam prom_inst_1.INIT_RAM_1B = 256'hD1F63DEAFA383B1D55EC77878B81CFEBEAF71FBFFFF3EE01D3BBEFFBBB65F8D2;
defparam prom_inst_1.INIT_RAM_1C = 256'h3D2BC72C3F22D6077790F1CFFFCCFFD065FBFF1FEECFC3B8FF8FF884EF4653BD;
defparam prom_inst_1.INIT_RAM_1D = 256'hFECAF2BA1F1BFA3737BDFDC8C3798576BDBFE7FFFE0EEEEFD4813C721EDAEF7D;
defparam prom_inst_1.INIT_RAM_1E = 256'hC0000330F403BC7E0C36FCA022B2EEE3BB6B2E03C23C70C13EBCC181AC48015B;
defparam prom_inst_1.INIT_RAM_1F = 256'h0C0C0EEB23CE34D30C34C00035D48022BB30440AF7E8C110AECCE0B860C38438;
defparam prom_inst_1.INIT_RAM_20 = 256'hA2D308031318C66000CE09F839C848AF8AC82EBFAF0AC433078B5CC281420AC8;
defparam prom_inst_1.INIT_RAM_21 = 256'h208C7CB9FA7F1C0AC8187ACC31ACC39124E20CFAD3933084A38F0BEE734806B3;
defparam prom_inst_1.INIT_RAM_22 = 256'hE812F22318EE327DAA20B20F18FF0E8FCAF8ACC00B002E8104EA302C8463CE28;
defparam prom_inst_1.INIT_RAM_23 = 256'h8F822F9E9E2BF67E7D86B13132F7810440000FC03F00FC4FF83A3E1B0004FF82;
defparam prom_inst_1.INIT_RAM_24 = 256'hCA32102D03B00F4C00A08C20310EB4103BCE732AEEB3AECEBCCAF1BC46B3BCEB;
defparam prom_inst_1.INIT_RAM_25 = 256'h80F33C12010032010424FC232304EC89E4F22CBAB02488AAAD48728CEB284A3B;
defparam prom_inst_1.INIT_RAM_26 = 256'hD0CCE31EC80C331C84312E111E28CBC000DCA7B03C3C3838360C00208038800F;
defparam prom_inst_1.INIT_RAM_27 = 256'h63CA00CC591CC0C3CB2CB91CC02CB2C412C3B38CBB000343722CB2CB2E4A30CC;
defparam prom_inst_1.INIT_RAM_28 = 256'h3E7C331CE4830D44330CC43F0A2ECA3D830D844B12C4F03C0A2CCA3D8DDEAD19;
defparam prom_inst_1.INIT_RAM_29 = 256'h9A86A1B00093139041F85C5D51DB6D79EF9EDA6CEC6CCE6C6C6C4E4C4E01CE5D;
defparam prom_inst_1.INIT_RAM_2A = 256'h31C59D2BA43036BDAB7BDE57BB4B8E60259025AE50A01A6163065A6126F39113;
defparam prom_inst_1.INIT_RAM_2B = 256'hFAA984E6E00474200034AC62C62F4990C0CE61984BE9631AD64D198F195C4052;
defparam prom_inst_1.INIT_RAM_2C = 256'h087E4975F07FCBC0CC147AB03C2E7F8D3C7EEEEF227F4B1CE8AEA67F0B2E17E6;
defparam prom_inst_1.INIT_RAM_2D = 256'h7641F41F86EB13E38F25D3E326CEC6CCFC01FE389104FC71E9BCF1FBC92C593A;
defparam prom_inst_1.INIT_RAM_2E = 256'h3844E11C81F579F94631CD87D34F8DFF3453E7F8D1371C9A82AAD358F1F93818;
defparam prom_inst_1.INIT_RAM_2F = 256'h7186CD5BE63073C798F873E61D3C0000344D6355388561352090D1E666307369;
defparam prom_inst_1.INIT_RAM_30 = 256'h0932CB0B16134C00AC04F08300180E44EC96CDC9206E67C98AE30003C4E4F002;
defparam prom_inst_1.INIT_RAM_31 = 256'h0000000000000000000000000000000000020585D3002805D300243A227C98AB;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[29:0],dout[5:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 2;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'hCEB2900E903B130B2AA0A92F8F037F385BF188CE23CAAAA00E0CEC2200333FC0;
defparam prom_inst_2.INIT_RAM_01 = 256'hC4301CC720C0720C4302CE00E084080323E007F3CAC8CF09300AC8EC8D380C18;
defparam prom_inst_2.INIT_RAM_02 = 256'h303333A3088FCB0438210004805FC48457F8484D3C4210204809FC84805FC411;
defparam prom_inst_2.INIT_RAM_03 = 256'h8C3CB00030C2CC4300FFCCCFCC400B3108CF03088788C3CE001100100C832033;
defparam prom_inst_2.INIT_RAM_04 = 256'h804423CF3130032C33733330C3C8CAE00334300820EB33040CF3CC4C818CE80E;
defparam prom_inst_2.INIT_RAM_05 = 256'hC886CFDB2CF04CC00CC30B8800CA123BC62C50BE03A8E310EA3BBCA084CAA280;
defparam prom_inst_2.INIT_RAM_06 = 256'hB34100001813C94F2020CC3CB00013101809002003BE10C020CF3CB02C80C8F2;
defparam prom_inst_2.INIT_RAM_07 = 256'hE33C001C400CCB01CCC93074103C18F0113FC0730F8CBCFF4B300C0C853CC3B4;
defparam prom_inst_2.INIT_RAM_08 = 256'h018000E28CF3C8300CC8A30C20414E32303308208CF3C4F0488CC34C34C32A30;
defparam prom_inst_2.INIT_RAM_09 = 256'h0040000000BFFFFF00EFEABA00BEAFBE00EABEBF00042450381059E0000F2687;
defparam prom_inst_2.INIT_RAM_0A = 256'h0400000000400000004001100000000000000500040504100110000000000000;
defparam prom_inst_2.INIT_RAM_0B = 256'h0004000001100040000000001014051400010550041501400401140400000554;
defparam prom_inst_2.INIT_RAM_0C = 256'h0554155515551555155505000000155505541555155510010554155515500554;
defparam prom_inst_2.INIT_RAM_0D = 256'h4000001000000004000014010005140505550015055500010414155505541555;
defparam prom_inst_2.INIT_RAM_0E = 256'h0554155515551000155515551555140515550154155514000555155515541555;
defparam prom_inst_2.INIT_RAM_0F = 256'hFFFF005505550404155504041555155515551515101500050554155510141555;
defparam prom_inst_2.INIT_RAM_10 = 256'h1C4711CC730C8320C8320000418C00AF8A0BF10000010400C10410410400C30C;
defparam prom_inst_2.INIT_RAM_11 = 256'h0A108184206104000014A0A0A0865B6C82188880CC400C8730C8330C4330C031;
defparam prom_inst_2.INIT_RAM_12 = 256'h6C718AAC22ACA81A18768C12EC410C4105387FC6A13C8F22108204C104C42202;
defparam prom_inst_2.INIT_RAM_13 = 256'h310E10210138400730C00733CF8C41421023CCF10F13C1A801843C4F30410434;
defparam prom_inst_2.INIT_RAM_14 = 256'h0E233CA10E30808428828418808428020850802A0A0A30E30CC0184C0D01384C;
defparam prom_inst_2.INIT_RAM_15 = 256'h320081313131313912C000002104F38C047012C03CCF0E123CE101384086A006;
defparam prom_inst_2.INIT_RAM_16 = 256'h4830F083822F0288C400003000213C0F12000C71081C4300CC004043C304C4C6;
defparam prom_inst_2.INIT_RAM_17 = 256'h00C484700320E1080003A200E0F18C28280F0A01C3002208283E4EC20F200218;
defparam prom_inst_2.INIT_RAM_18 = 256'hA000204C4C00820000100204C808C30820CC8231208000043208F02043128493;
defparam prom_inst_2.INIT_RAM_19 = 256'h0A82102102100C2080003202080201F06F2330C420C8F2080080F208C3002210;
defparam prom_inst_2.INIT_RAM_1A = 256'hC4F80320C03000000026CC0054A8D7345314D81F16C0422A8822C302030A0802;
defparam prom_inst_2.INIT_RAM_1B = 256'h14C53607C5B0C8300020C040888B100301C43081320030931000030008420413;
defparam prom_inst_2.INIT_RAM_1C = 256'h3A03FF303F3108C4C8307307108000320208134200204800CC41023700DCDC03;
defparam prom_inst_2.INIT_RAM_1D = 256'hCF01C03C30DF3CC808023026CC3F3001321334C00440000204033CF3120633A0;
defparam prom_inst_2.INIT_RAM_1E = 256'hAAAAA83AAFBAEBEA2EEEAA82AAE8000004040F90E380081B43C01B5B73114867;
defparam prom_inst_2.INIT_RAM_1F = 256'h0D4C4E08830C30C30C30C2AAAABEBEAAE03BBAABBAA0EEEABBAE82EA82EAAAE8;
defparam prom_inst_2.INIT_RAM_20 = 256'hA61990A63B72DCD5258D63D973D69611A116700C11211E508DAC610F23012112;
defparam prom_inst_2.INIT_RAM_21 = 256'h7A194181384E4DC11661B021000210070AC018F12758458D4B56403B54110008;
defparam prom_inst_2.INIT_RAM_22 = 256'h0449471071D652048549442B50F69D41911A11201C427045942112614D0BE684;
defparam prom_inst_2.INIT_RAM_23 = 256'h01A714131300804C4E81C4B99949A01CA00903E40F903E721A75065C555721A6;
defparam prom_inst_2.INIT_RAM_24 = 256'hD83500849C52712482850151B50D055270DCF7200008001CBDC00B0CDC751D43;
defparam prom_inst_2.INIT_RAM_25 = 256'h33370C6071716140144200462050009802030000478DC19AA05B76DD736F5CB2;
defparam prom_inst_2.INIT_RAM_26 = 256'hE50103500A0D4071410470143E7D1028141DC33D0D0D0D0D0F40108CC102033F;
defparam prom_inst_2.INIT_RAM_27 = 256'h036D840D1351026FD0410351024104142414C50D48042394C72D041040DC3500;
defparam prom_inst_2.INIT_RAM_28 = 256'h087C3B0EDE1041410B42C10F91511162104182D0B400F90C515111620A52CF15;
defparam prom_inst_2.INIT_RAM_29 = 256'h164591CA95001138E14372525710410030D34C0E0E4E4CCECECECC2264429041;
defparam prom_inst_2.INIT_RAM_2A = 256'hB5C44DC3C509363D0B62DCD0019F6D724F5C8F3C63C91450509D14F009E73BBB;
defparam prom_inst_2.INIT_RAM_2B = 256'h04E49415004D4512EED63E53E53D635C24ED735852D35098D02C1D4B43415161;
defparam prom_inst_2.INIT_RAM_2C = 256'h1896550612416248659AF7D735D3711412A2222496711514D5D2967115123615;
defparam prom_inst_2.INIT_RAM_2D = 256'hDB414514252899597D76105971E1E5E5D601059139C416535E165AA1694E3D95;
defparam prom_inst_2.INIT_RAM_2E = 256'h94121150190942F3E50BA25715B9790599413416454734D146AA6E55F2A5C490;
defparam prom_inst_2.INIT_RAM_2F = 256'h43572771F71351CF9CB562D43CB49EEEDA705700B419D1866554554D4D534151;
defparam prom_inst_2.INIT_RAM_30 = 256'hA94A69A5011C268215871A49A0864F8526A420685D410F6A3C5EEEED67161A08;
defparam prom_inst_2.INIT_RAM_31 = 256'h000000000000000000000000000000000001004709A0844709A0993C94F6A3C9;

pROM prom_inst_3 (
    .DO({prom_inst_3_dout_w[29:0],dout[7:6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .AD({ad[12:0],gw_gnd})
);

defparam prom_inst_3.READ_MODE = 1'b0;
defparam prom_inst_3.BIT_WIDTH = 2;
defparam prom_inst_3.RESET_MODE = "SYNC";
defparam prom_inst_3.INIT_RAM_00 = 256'h7010402C6C3D604D301AC3B1EC3EEDB3F37FFFECCE4FFFF02CC2C00F0DF08733;
defparam prom_inst_3.INIT_RAM_01 = 256'hF73DCF33CCF33CCF33CCECDEC03333DD0B13FFDE787BAC7FFEC0774777B0370F;
defparam prom_inst_3.INIT_RAM_02 = 256'h0EF00B3F3BB5EC7BB00CC0374F7F774F736374F33770DCCF74F3F4374F3B77DC;
defparam prom_inst_3.INIT_RAM_03 = 256'h7BB2CFCFF3F3C37EF3FFC3FFC37DCF0DFFACEF3FB4FF7B13EFEC3FEC7FCDCEF0;
defparam prom_inst_3.INIT_RAM_04 = 256'h73B0DFCF0DF37BB3F08F08EF7B3F71AC01CC30F7CFF30EF333F3C37C730CC73C;
defparam prom_inst_3.INIT_RAM_05 = 256'h37ECACF3B2CCEF7DEFBEECB7EC2CDFB1FFFFB2CFFB02CED2C0B032CFFB2CFB3F;
defparam prom_inst_3.INIT_RAM_06 = 256'hF043C000CFF7F3DFCC0EFFB2CFDCEF03FFFFFFEFFB3CDEFFEF33B2CBB333F73B;
defparam prom_inst_3.INIT_RAM_07 = 256'h1DF003FFF3BC0DEDC0CD107FEDB3FACEC0B33B3EECBBF7B94F0FDBB8F7BC11D4;
defparam prom_inst_3.INIT_RAM_08 = 256'h00BF33FB37CB373CCF3ECFF3CECE34CCCF35F3CC079E73CF333770770770B1DC;
defparam prom_inst_3.INIT_RAM_09 = 256'h002A00000000000000155555001555550041555500020002015550000FEC0438;
defparam prom_inst_3.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam prom_inst_3.INIT_RAM_10 = 256'hDFB7FDF37DDFB7EDF37FF7DF3D33DE872CC1CFFF0FBEFB0F7DF3EF7CFFFF7CF3;
defparam prom_inst_3.INIT_RAM_11 = 256'hE8CF7A33DE8CFF3CF0F28E8E8F7311473DCFB3FCD73EDF77CDF37EDF37EDF77E;
defparam prom_inst_3.INIT_RAM_12 = 256'h868A28000A3E8FA3A310F3DF477DF37D28028C68FDE739FCCF3FFB7CFB73C47D;
defparam prom_inst_3.INIT_RAM_13 = 256'hCCE8CF8CECA3F3FFDC03FFDF2C833B2CCF8B3B9FECFE7A17BFF3B339CF7DF702;
defparam prom_inst_3.INIT_RAM_14 = 256'hECF00C3CF8DF7A33E37B33E37A33D37DF35A3BB3A3A1DC1DC3FCC33BF86CA33A;
defparam prom_inst_3.INIT_RAM_15 = 256'hFCCF3FDFDFDFDFDFFF33CF3FCFFF9A3B3FC0FF33B3B9C0EC368CECA33E285EFF;
defparam prom_inst_3.INIT_RAM_16 = 256'hBF3A13730DCD093F73FF0FD3F0CCE779CCFF768CF3A373DCF35F33F0CDFF7F68;
defparam prom_inst_3.INIT_RAM_17 = 256'hDFF3F44A68EF4FC334E80DFF0A3FFB0E8339A35A28DFCFA28E87F468A1FD68FF;
defparam prom_inst_3.INIT_RAM_18 = 256'h4FBFCFB7B7DC3CFDF7ECFCFB77F78CC3CC733CDCCF3F7DFBDDF39FCFBDECFBFF;
defparam prom_inst_3.INIT_RAM_19 = 256'hA168CE8CE8CCA093BDF7EC3CF3FC3F7FCD6EEA10DFF30EF3EFB67EF3D903DFCF;
defparam prom_inst_3.INIT_RAM_1A = 256'h7793F5ECFB30000000DCF3A35E4F33CF37CDDF73CCF3318033CCF300E8A3A168;
defparam prom_inst_3.INIT_RAM_1B = 256'hCDF377CCF73FBFCD00FF3FFFB3B1FFF3FCF7CF3EDDF7CFFDDFF0FD3F037CF7DE;
defparam prom_inst_3.INIT_RAM_1C = 256'hF1DFFF0EFF0DFFF7F7CF3CF3DF3DF7CC3CF3ED0DFFC333FCD77CF4CFFDCF3FF7;
defparam prom_inst_3.INIT_RAM_1D = 256'hECCCF337CFFFB3FFFF0FD3FCF737CCFF33DED7B007FFDFDEFF7CFCF0DDEC331E;
defparam prom_inst_3.INIT_RAM_1E = 256'h0000000155155555005554005553FC3FF0F0CDFEC33333010B330101102083FE;
defparam prom_inst_3.INIT_RAM_1F = 256'h0141405100410410410410000554545550015505555005545555401540055454;
defparam prom_inst_3.INIT_RAM_20 = 256'hFED1370DE1DCF78DC378DE70DE7CF0CF0CFCFF30CF0CF8CC0300FF3900030CF8;
defparam prom_inst_3.INIT_RAM_21 = 256'hE3FBDFBCD33537FCFCFCDCC3B0CC3B0FCF403BFCFFF3F3BBB30C0040555FB331;
defparam prom_inst_3.INIT_RAM_22 = 256'hF3F33DFBDDCC345D33F37DC3DCDC3FCF0CF0CF8CFFCFFF3F3EFCF0EF3B334C33;
defparam prom_inst_3.INIT_RAM_23 = 256'hCF0FF3CDCDF30F3737C659111F3F003FC0C3F74FDD3F74CC30FF3C33F3BCC30E;
defparam prom_inst_3.INIT_RAM_24 = 256'hFB30003D37F4DF4D00FF70DC0DCC0CCCFCFF9FCCC330CC3F37FCD1CC333CDF33;
defparam prom_inst_3.INIT_RAM_25 = 256'hF00FC0C1C1C1C1C178545054005414115450400F3E3373B004FB3ECFB3ECF73C;
defparam prom_inst_3.INIT_RAM_26 = 256'hFCD3B3CD08CF34FF7330FF3DE4DA73428CE3387F373737373DCC003C033FC30C;
defparam prom_inst_3.INIT_RAM_27 = 256'h33D3FDCCFECD00D333CF3ECD00CF3CFF7CF34ECF34400FF34DEF3CF3CFB73CD3;
defparam prom_inst_3.INIT_RAM_28 = 256'hBB7771DC70F3CF7331CC433CF3CD33FFF3CF30731CC3FF7C33CD33FFC1587007;
defparam prom_inst_3.INIT_RAM_29 = 256'hE0380FF000CCCCC30FFFEFEFFF3FFFFD965967646464676464646744470048EF;
defparam prom_inst_3.INIT_RAM_2A = 256'h037ECFB37DC0EDCFB3DCF7B70FF7DCCC393332E7CE40E3CCCC0433903659E221;
defparam prom_inst_3.INIT_RAM_2B = 256'hDF3F3CFFD0337CF04470E4FE4FE70E3B0380EE37DCCEEC3BBB0137B30EDCDCDC;
defparam prom_inst_3.INIT_RAM_2C = 256'h0030EFFEF0EF0EC04C343C30CC30DF0C3058888C30DF0C330C30F0DF0C30CDFF;
defparam prom_inst_3.INIT_RAM_2D = 256'hB0DFBCFBFFC111C3030DFFC30646464670033C30CFBCF0FEC3F0C16F0FB23513;
defparam prom_inst_3.INIT_RAM_2E = 256'h10044037FF7FDFDCBDC283FFFF0B0B3C30DF0CF0C3BCEC3CC000C2CCC06FFC33;
defparam prom_inst_3.INIT_RAM_2F = 256'hEE3CC4FDDFF0FDC13F30FCCFE51C344470DFFC00D00FBF3FF03B73B8F830EDCD;
defparam prom_inst_3.INIT_RAM_30 = 256'h0F3FC30CC3FFFC00F3FFF0C3003DCDFCFC3CF5C3F7CF79C3E7C244470DFCF003;
defparam prom_inst_3.INIT_RAM_31 = 256'h000000000000000000000000000000000003B0FFFF003EFFFF003B37FB9C3E7F;

endmodule //t20k_rom
