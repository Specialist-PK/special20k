//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.10.03 (64-bit)
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Tue Nov 26 22:45:02 2024

module t20k_rom (dout, clk, oce, ce, reset, ad);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input [12:0] ad;

wire lut_f_0;
wire lut_f_1;
wire [27:0] prom_inst_0_dout_w;
wire [3:0] prom_inst_0_dout;
wire [27:0] prom_inst_1_dout_w;
wire [7:4] prom_inst_1_dout;
wire [23:0] prom_inst_2_dout_w;
wire [7:0] prom_inst_2_dout;
wire dff_q_0;
wire gw_gnd;

assign gw_gnd = 1'b0;

LUT2 lut_inst_0 (
  .F(lut_f_0),
  .I0(ce),
  .I1(ad[12])
);
defparam lut_inst_0.INIT = 4'h2;
LUT3 lut_inst_1 (
  .F(lut_f_1),
  .I0(ce),
  .I1(ad[11]),
  .I2(ad[12])
);
defparam lut_inst_1.INIT = 8'h20;
pROM prom_inst_0 (
    .DO({prom_inst_0_dout_w[27:0],prom_inst_0_dout[3:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_0.READ_MODE = 1'b0;
defparam prom_inst_0.BIT_WIDTH = 4;
defparam prom_inst_0.RESET_MODE = "SYNC";
defparam prom_inst_0.INIT_RAM_00 = 256'h4A1E955559119F6A02218B55555555301FAA001F6290015500443F322EFF1033;
defparam prom_inst_0.INIT_RAM_01 = 256'hB2D99906FA086F82706FFC6CF15EF36C0B999F5F7A06F929BFD236022EECFCA0;
defparam prom_inst_0.INIT_RAM_02 = 256'h06FC2FA60425ED91E96F90F27FAAF911110C25D5713DB4713DA1F8A860625350;
defparam prom_inst_0.INIT_RAM_03 = 256'hE1AACE17AAE1BA9E1DA8E17A8E18ADE13AAE17A0EFCA013FC208100D02DD0A3C;
defparam prom_inst_0.INIT_RAM_04 = 256'hDA1EDD61D373619A2EC1D30617302DD1D3FA61125ED061D3736132EEC1D317AF;
defparam prom_inst_0.INIT_RAM_05 = 256'hAE1FDF32BEF1A55509E03A9FEF9AF0E3FC208100D00001D3FA61D25ED1D3FA61;
defparam prom_inst_0.INIT_RAM_06 = 256'hD12A7F4A23DF655133FE59110DF120E5273110D56599102559111016251FDF32;
defparam prom_inst_0.INIT_RAM_07 = 256'hF153F42FCA1A251A3F612226F1A24D153252FE06F2A1F2FEF0A2AD2BA26F1A24;
defparam prom_inst_0.INIT_RAM_08 = 256'h777927AFCDE0920426D976FF1A1532225252FE36F1A24DF692AA9CBEFE7283F6;
defparam prom_inst_0.INIT_RAM_09 = 256'hB2D10D56292FE36F1A24DFE31A0EFFA59F321E9F322E15310DF42911E46F5067;
defparam prom_inst_0.INIT_RAM_0A = 256'h5555911214FFAA5591FC2BBFCA2CDFEFC233FCA4BF6FB159121C5FB159FDA912;
defparam prom_inst_0.INIT_RAM_0B = 256'hA37A9FFA7F4A581EFF2F023A21E10D3EA0E20D11DFA2F20D23D16FB1003BFCA9;
defparam prom_inst_0.INIT_RAM_0C = 256'h11128D5552831BD283FA2FF1372CE28310D31AAEF42FC206FCA33209130AAEFC;
defparam prom_inst_0.INIT_RAM_0D = 256'h6F1A70E55000000090E2820E190680E13B30010BE203F0AFF291332D10DF60E9;
defparam prom_inst_0.INIT_RAM_0E = 256'h2596F32FE3229E3C3F32F3226E93E27AF16F1A39DF137AB164AA0EF1AF7F69F1;
defparam prom_inst_0.INIT_RAM_0F = 256'hEF37DFE00009111362D48DF321EB48DFF32E61677A8E75551037FFA9119F3A32;
defparam prom_inst_0.INIT_RAM_10 = 256'h07D80EFE94D247D332E9BD0AC463FE9442347D737D8E737D8EF37D8EF32737D8;
defparam prom_inst_0.INIT_RAM_11 = 256'h000802800002C9F1A393FEFF24FAAE80ADE37D9F3A39D48D4DDFF14414314833;
defparam prom_inst_0.INIT_RAM_12 = 256'h0000FFC02849D3E10000DA8080B9A9C10F0D127F200FC800003C3FEA00F0016A;
defparam prom_inst_0.INIT_RAM_13 = 256'h0000FCBA765432100000D0987654321B0000A8ADB7E5B53A0000EC64CF201796;
defparam prom_inst_0.INIT_RAM_14 = 256'h000042660D25CAA40338429804E5E4F40AAFAFAA00000AAA0404444400000000;
defparam prom_inst_0.INIT_RAM_15 = 256'h000842100CC000000000F000084CC0000044F4400045E5400842224802488842;
defparam prom_inst_0.INIT_RAM_16 = 256'h0888421F0E11E0870E111E0F022F2A620E11621F0F08611E0E4444C40E19531E;
defparam prom_inst_0.INIT_RAM_17 = 256'h0404211E08421248000F0F0002480842084CC0CC0CC00CC00C21F11E0E11E11E;
defparam prom_inst_0.INIT_RAM_18 = 256'h0F13001E0000E00F0F00E00F0E99999E0E10001E0E11E11E011F11A40E07531E;
defparam prom_inst_0.INIT_RAM_19 = 256'h0E11111E01135911011155B10F100000012484210E1111110E44444E0111F111;
defparam prom_inst_0.INIT_RAM_1A = 256'h0A555111044AA1110E1111110444444F0E11E01E0124E11E0D25111E0000E11E;
defparam prom_inst_0.INIT_RAM_1B = 256'hF0000000000001A40E22222E001248000E88888E0F08E21F04444A11011A4A11;
defparam prom_inst_0.INIT_RAM_1C = 256'h0000001F044F55F40F02E20F01FAAAA601F222220E11E00F011F111E0255D552;
defparam prom_inst_0.INIT_RAM_1D = 256'h0E51115E0111F111011155B109999997013484310119531501195311011A4A11;
defparam prom_inst_0.INIT_RAM_1E = 256'h0E11E11E0155E5510084A1110E44445F0E10001E0000E11E0195F11F0111111F;
defparam prom_inst_0.INIT_RAM_1F = 256'hFFFFFFFF0111F11101F555550E11711E0F5555510E11611E095591110E11E000;
defparam prom_inst_0.INIT_RAM_20 = 256'h1F12801FF18238E3009C939B3903009AC3EC3ED3ED3EC3BA3303E83373373863;
defparam prom_inst_0.INIT_RAM_21 = 256'hA2E9BA7E86A8ECBA4ECAABECDACED5ADEEFA4EC1DF3DD9DEDDF218638BDFB2EF;
defparam prom_inst_0.INIT_RAM_22 = 256'h9DCCD958D33E5D80EFEE43A0AFEB1A3EC2A6E94A7E92A9EC6AEE89A8EC6A3E90;
defparam prom_inst_0.INIT_RAM_23 = 256'hDF5A98DCCDF7A98DCCDFDA98D8E2D193D54EF61F419FBA9FB29CCD9137FAFFBE;
defparam prom_inst_0.INIT_RAM_24 = 256'h1FA1081F92F6EF72B591A7A9E27B9B13EDDE9D5B9EDD9198DEDD898D5BEB69CC;
defparam prom_inst_0.INIT_RAM_25 = 256'hA17F9AF7AF52339001F3215F1215FF2BFD292E33986397D11B098D98D369AD9D;
defparam prom_inst_0.INIT_RAM_26 = 256'hEDDF11FF29AA7DA83FE2A8A791F3290C9D555AA3FF2AAA7D86398D98D9AD081F;
defparam prom_inst_0.INIT_RAM_27 = 256'h1AEDDF01EDDFE144DF01F019B2D9B29E37D8E2E9B29E37DFEF32F06BADF01F11;
defparam prom_inst_0.INIT_RAM_28 = 256'h247D09FAAC9DF3ABFC2BFA2737D8EF37D8E39DAB333AAA79B29AEF11F01AAA7F;
defparam prom_inst_0.INIT_RAM_29 = 256'h9FCA91C6D6F315EDDFC1A23CCDFCAEDDF91CCDF3AEDDF61CCDFAAEDDF01F3DAC;
defparam prom_inst_0.INIT_RAM_2A = 256'hD30D9E3E30D6EBEDFE2A0A79106BAD23DEEF01BADF01F01EDDF11F3290C9D555;
defparam prom_inst_0.INIT_RAM_2B = 256'hA233B0A47D30DE30DA30DB30DC30DD1130D6EBEDBEDBEDA63330DA2A7EF01AA2;
defparam prom_inst_0.INIT_RAM_2C = 256'hBC331E8DF57F5ABCA47DF52BFADEB0A8E37DD49B02D30D0EFEA2330DC30DDF3A;
defparam prom_inst_0.INIT_RAM_2D = 256'h9A111EF929DB82DE3CBF2CEE0EF015597BC31E8D8EE8DFEE8D8E5BBCA9DBA28C;
defparam prom_inst_0.INIT_RAM_2E = 256'hE23C729EFEA5E7F02F9AEDD847D1FE2FA15FA29111133FC1FB2DC9D4DF7A555B;
defparam prom_inst_0.INIT_RAM_2F = 256'hF3DB62DE5DFEFD007F9A8DDF41BE253CCD746F9ABBCCDBE2DBF9A5555B32531F;
defparam prom_inst_0.INIT_RAM_30 = 256'h47D2EC233847D1C633847D1F3DEDDEDD5ECCDCAA9E91E9DEDD5EBD331BD31111;
defparam prom_inst_0.INIT_RAM_31 = 256'h015C9D91E9DEDDDEDDC5C6333847D1F3DEDDEDDA51E9DEDDECCD5C3AEACB3338;
defparam prom_inst_0.INIT_RAM_32 = 256'hA0E9F1CCA7F5AE06CCD9193933C9247DCC3C0D7E81CBA47D5F1E0019CCD1EDDF;
defparam prom_inst_0.INIT_RAM_33 = 256'hF7209F52D0DF32D0DF12D0D3F02AF01CD3F3DEDDC2235847DE9DE8DEEC9AFEC7;
defparam prom_inst_0.INIT_RAM_34 = 256'h427EE4A1EF6D4AAEE4A0E93D333F59999DBDD9ACE8DEA0019F0AF1ABF3A4DF5A;
defparam prom_inst_0.INIT_RAM_35 = 256'hDD428C3E8DF7D0ADED7A8E00000000000000D3A1E37DF0154D5F01590606976E;
defparam prom_inst_0.INIT_RAM_36 = 256'hD9AAEE6D37DE9DEDDECCDF3DFBD91117D43E8D8EE8DFEE8D8EBD4A47DE93D429;
defparam prom_inst_0.INIT_RAM_37 = 256'hE427EE4A1EF6E9AAEE9A0E910DAD37D77777DAD37D5D935D83BD8337D1DDDA8E;
defparam prom_inst_0.INIT_RAM_38 = 256'h5847DE9DEDDE06CCD9E8D0EED33E8D80EFEE93EDDF919061E8DF5069761E8DF5;
defparam prom_inst_0.INIT_RAM_39 = 256'h3FE728AFE06F2AE22FEF0A2AD559124D5E5D8630FE37D0FEECDEF3F3DEDDE423;
defparam prom_inst_0.INIT_RAM_3A = 256'hAEF69FECDB7ECDFFFFF911E8DBE8DAEDD55283252FE36F1A24D9E7A9CBEF6FE5;
defparam prom_inst_0.INIT_RAM_3B = 256'hEFDAF2AAEF2AAE9907DE148EFCA91E5D1E5D8EE5DFE5E0A0E10C7E9590676E5A;
defparam prom_inst_0.INIT_RAM_3C = 256'h8D9E59AE0AE9111FC2081FD25F02D3370EFAAFF2D337A337A8E060A10015558E;
defparam prom_inst_0.INIT_RAM_3D = 256'hE0000000000D0D01DD53011E8CF24EFB00F02F49EFD0AA011B29BF09E8DAE91E;
defparam prom_inst_0.INIT_RAM_3E = 256'hBFAD0D03524100A9EE5EFBA0D0352410A9E8C1E1EA00ACA16A00F01CA1601D90;
defparam prom_inst_0.INIT_RAM_3F = 256'h00D030D300D9C88D0A0DC0D80D50D40D30D20D60D10000000E54F77092001B29;

pROM prom_inst_1 (
    .DO({prom_inst_1_dout_w[27:0],prom_inst_1_dout[7:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_0),
    .RESET(reset),
    .AD({ad[11:0],gw_gnd,gw_gnd})
);

defparam prom_inst_1.READ_MODE = 1'b0;
defparam prom_inst_1.BIT_WIDTH = 4;
defparam prom_inst_1.RESET_MODE = "SYNC";
defparam prom_inst_1.INIT_RAM_00 = 256'hDD2F7FCDECECF8F2C2CB70EEEEEEEE0008F2C038F23002CE00C4CF03837F3C0C;
defparam prom_inst_1.INIT_RAM_01 = 256'h7C322702610008F269C00FE7490340E70E222688E22D8E37E8F30CCBDBF78F2C;
defparam prom_inst_1.INIT_RAM_02 = 256'h028F360CCCDFF7CB7CA27CACB8F34CEDCFC8C0227C6C727C6C7D8F200C7C01EC;
defparam prom_inst_1.INIT_RAM_03 = 256'hFC5C0FC4C1FC3C1FC2C0FC0C1FC2C0FC1C0FC0C2F8F2C4C8F2002C1C0C2CC4C7;
defparam prom_inst_1.INIT_RAM_04 = 256'h5D1F7B2C5C60DC3D0F7C5C02C5C0C2CC5C60CC2DFF702C5C60CC1DBF7C5CC5C1;
defparam prom_inst_1.INIT_RAM_05 = 256'h03C8CF03038F2ECF0CACAC77F8E34C9C8F2002C1C0000C5C60CC5DFF7C5C60DC;
defparam prom_inst_1.INIT_RAM_06 = 256'hCCECB8F3C8CF0CECAC53ECEC7C8F343EC8CCC9C10CCCC9C04CFCE0C7C2C8CF03;
defparam prom_inst_1.INIT_RAM_07 = 256'h6CBC8F38E3CCC0CCCF0CFC0EF03C5CCBCC0CFFFFF03CFCFFF03C5CC4C0EF03C5;
defparam prom_inst_1.INIT_RAM_08 = 256'h0007C3D00F00CC6CC2CCFE2F03CBCC1C0C3CFF0FF03C5CF06C0D20F0F26C0CF2;
defparam prom_inst_1.INIT_RAM_09 = 256'h6C0C9C10C6CFF0FF03C5CF0C4C8F8E3CCF0393CF0383CBCC7C8F3CEC7C26BAC0;
defparam prom_inst_1.INIT_RAM_0A = 256'hFCDECEFC9D08E3FECC8F2228F2CBC508F2228F232F38E2CCEC9C38E2EE8E2CCC;
defparam prom_inst_1.INIT_RAM_0B = 256'h3C6CE8D2B8F3FD2F8E38F3C0D8FC7CC4C8FCBCCBC8E3AC6CC8C038E2C5CE8F27;
defparam prom_inst_1.INIT_RAM_0C = 256'hCDECCCEDCCCCCACCCC8F2FF2C5C8FCCCCACC3C3F8F38E38C8E3C2C0CFC6C3F8E;
defparam prom_inst_1.INIT_RAM_0D = 256'hEF03500DC0000000C1ECCD4FFC2DD4FFC2C002C8FCFC8F38E3CCC4C0C9CF010C;
defparam prom_inst_1.INIT_RAM_0E = 256'hC1018F3F3C8C1FCBC8F3ACBCEF7CBFB750EF03CCC4BC8CB0EC5D8FF03407E750;
defparam prom_inst_1.INIT_RAM_0F = 256'h36C7CF30000CCDFCDC0C8CF030E7C8C5F030F0E507005FDCC9C48F3CCDA8F3C8;
defparam prom_inst_1.INIT_RAM_10 = 256'hC3CC0F47CC2CC2C0207CB7CB7C1CF3CC1C2C2C7C7C035C7C035C7C038E26C7C0;
defparam prom_inst_1.INIT_RAM_11 = 256'h0001ACCC0C0CFE8E2C7CF38F3C6C0FC0C0FC3CE8E2CFCC3CC2C8D0C91C72C3C2;
defparam prom_inst_1.INIT_RAM_12 = 256'h00007226677667770000001802101108032445445521320000CCC8F302522C93;
defparam prom_inst_1.INIT_RAM_13 = 256'h0000188800000000000023333333333300003677766667660000277666776776;
defparam prom_inst_1.INIT_RAM_14 = 256'h0000000000110000001000110010010000010100000000000000000000000000;
defparam prom_inst_1.INIT_RAM_15 = 256'h0010000000000000000010000000000000001000000101000000000000000000;
defparam prom_inst_1.INIT_RAM_16 = 256'h0000000100111100001001110001100000100001011000100000000000111110;
defparam prom_inst_1.INIT_RAM_17 = 256'h0000001000000000000101000000100000000000000000000100011000110110;
defparam prom_inst_1.INIT_RAM_18 = 256'h0011111001111111011111110100000100111110011111110111110000111110;
defparam prom_inst_1.INIT_RAM_19 = 256'h0011111001111111011111110111111101111111001100000000000001111111;
defparam prom_inst_1.INIT_RAM_1A = 256'h0011111100000111001111110000000100100110011111110011111001111111;
defparam prom_inst_1.INIT_RAM_1B = 256'h1000000000000100000000000000001000000000011000010000001101100011;
defparam prom_inst_1.INIT_RAM_1C = 256'h0111111100011110011111110110000000111111011111110111111001111111;
defparam prom_inst_1.INIT_RAM_1D = 256'h0011111001111111011111110100000001111111011111110111111101100011;
defparam prom_inst_1.INIT_RAM_1E = 256'h0111111101110111010001110000001100111110011111110100011001111111;
defparam prom_inst_1.INIT_RAM_1F = 256'h3333333300001111001111110010001001111111001000100111111101111111;
defparam prom_inst_1.INIT_RAM_20 = 256'h28E2C027F3CDCCCC00CC8CC9CC9C00CC7CC5CC1CC9CC5CC1CCDCCCCC7CC3CC3C;
defparam prom_inst_1.INIT_RAM_21 = 256'hC5FC9C5FCDC5FC3C5FC7C4FCAC4FCAC4FC2C4FCECC4CC4CC1CC52C3CC4C8A27F;
defparam prom_inst_1.INIT_RAM_22 = 256'h2CC6C1ECAC2CECC0F47C1CC8C4FC6C5FC3C4FC2C4FCBC4FC1C4FCBC4FC4C4FC9;
defparam prom_inst_1.INIT_RAM_23 = 256'hC8A2C1CC6C892C1CC6C892C1CCDC0CC0CC00CD18A2C8A2C8A2CC6C1E1527527C;
defparam prom_inst_1.INIT_RAM_24 = 256'h0891032893F37892EEC5CB7C2CB7CEC2C1CC2CCECC9C7CC1CC9C7C1CC2424CC6;
defparam prom_inst_1.INIT_RAM_25 = 256'h9278938928A22230028A2EF8A2EC892E892C1712EC3CC5CE727C5CC5CC3C5CC5;
defparam prom_inst_1.INIT_RAM_26 = 256'hC1CC828F3CBCB7CDC8F3CDCB7C89266C8CCDEC1C8F3C1CB7C3CC5CC5CC5C0318;
defparam prom_inst_1.INIT_RAM_27 = 256'hC3C1C8B2C1CC82C1C8C18B2CDC0CCCDFC7C0300CCCDFC7CF38F3A03C1C8D18C2;
defparam prom_inst_1.INIT_RAM_28 = 256'hCC2C55882C8C8E2E882E8826C7C036C7C03CFCC0C12C1CBCCCB148C18B2C1CB8;
defparam prom_inst_1.INIT_RAM_29 = 256'hC8F2CE0303F02EC1CCB2C7CC6C882C1CCA2C6C8E2C1CC92C6C882C1CC62C4CC6;
defparam prom_inst_1.INIT_RAM_2A = 256'h0CDCD300CDCE3C0C8F3CBCB7C032C9C20F78B2C1C8C18B2C1CC8289266C8CCDE;
defparam prom_inst_1.INIT_RAM_2B = 256'hCFC2C0CC2CCDC7CDC7CDC7CDC7CDC7EDCDCE3C0CC0CC0CCCC2CDCCDCB78B2CBC;
defparam prom_inst_1.INIT_RAM_2C = 256'hC1C2CCCC4C7893C1CC2C893C5C0FC4C0FC3C44CC1C0CDC03F0C7CCDC7CDC7892;
defparam prom_inst_1.INIT_RAM_2D = 256'h9CEC0F88370C6C0F20C6C2F700862CEC7C1CCCCC00CCC70CCC00C2C1CB7C4CB7;
defparam prom_inst_1.INIT_RAM_2E = 256'h822C0CB7882E44893883C4CCC2CE882882E8837EDC7278828837CEC44882CDEC;
defparam prom_inst_1.INIT_RAM_2F = 256'hC4CCFC1CEC5053884883CACC72CDC02C0C40C88322C6CCCC32883FCDECBC02E8;
defparam prom_inst_1.INIT_RAM_30 = 256'hC2C07C3C2CC2C7C1C2CC2CCC4CC4CC9CC7C6CC2CB7CCC2CC9CC7C9C2EC9CEDCF;
defparam prom_inst_1.INIT_RAM_31 = 256'h62CC8CCCC2CC9C7C9C7CC4C02CC2CCC4CC4CC9C0CCC2CC9C7C6CCC6CB0C3C02C;
defparam prom_inst_1.INIT_RAM_32 = 256'hD2F74ACBCB883410C6CCFC2C33CACC2CC8CCAC487FCACC2CF487000CC6CEC1CC;
defparam prom_inst_1.INIT_RAM_33 = 256'h88266882C1C882C1C882C1C08830860CACC4CC4CCBC20CC2CC2CCCC20CCD7FCC;
defparam prom_inst_1.INIT_RAM_34 = 256'h1D4FC1D4F5EC4D3FC1D2FC0C1C0682222C2CC2C2FC0F0002C883882E88244882;
defparam prom_inst_1.INIT_RAM_35 = 256'h7C5CB72CCC47CAC0FC8C0F00000000000000C6D2FC3C880C55D862EC3D1FC3DC;
defparam prom_inst_1.INIT_RAM_36 = 256'hCCC1FC5CC3CC2CC9C7C6CC4CC3CCEDC7C5CCCC00CCC70CCC002C5CC2CC5CC5CB;
defparam prom_inst_1.INIT_RAM_37 = 256'hC1D4FC1D4F5EC0D3FC5D2FCCBCECC3C40000CECC3CCCDCCCAC2CAC27CDCCCC0F;
defparam prom_inst_1.INIT_RAM_38 = 256'h0CC2CC2CC9C710C6CCCCC20C1C2CCCC0F47C5CC1CC42C3DFCCC4F1FC3DFCCC4F;
defparam prom_inst_1.INIT_RAM_39 = 256'hCF26C4CFFFFF03C8CFFF03C5CCECFC5CFC6CC3CC1FC3CC1FC5CC2CC4CC4CC3C2;
defparam prom_inst_1.INIT_RAM_3A = 256'h0F0EC5CBC75CBC00005CDCCCC4CCC4CACCDC4CC3CFF0FF03C5C6C8D20F0F26C8;
defparam prom_inst_1.INIT_RAM_3B = 256'hF8F3C0C1FC0C0F7CC3CCFDFF8F3CFCECCCEC00CEC70CCED2FC7C0F7FC3C0CCCD;
defparam prom_inst_1.INIT_RAM_3C = 256'hCC10CC10C0F7EDC8F20F2C0C0C2C0127108F3C0C0127112717030901902CDEDB;
defparam prom_inst_1.INIT_RAM_3D = 256'h2222222222200326667727667667766602327676666220026666762CCCC00CCC;
defparam prom_inst_1.INIT_RAM_3E = 256'h7600032767662267676666003276766267676676600236666002326666627660;
defparam prom_inst_1.INIT_RAM_3F = 256'h0035503450324424200340340340340340340340340222222266677267726666;

pROM prom_inst_2 (
    .DO({prom_inst_2_dout_w[23:0],prom_inst_2_dout[7:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(lut_f_1),
    .RESET(reset),
    .AD({ad[10:0],gw_gnd,gw_gnd,gw_gnd})
);

defparam prom_inst_2.READ_MODE = 1'b0;
defparam prom_inst_2.BIT_WIDTH = 8;
defparam prom_inst_2.RESET_MODE = "SYNC";
defparam prom_inst_2.INIT_RAM_00 = 256'h230036DE2A21380ED537CDD00CC2B0790B230036070001D90021C818CDD07E21;
defparam prom_inst_2.INIT_RAM_01 = 256'h7ED21F21E5D01821D1A7CDC809CD3E0EC818CDDD0021C818CDD1FB21D01DC20D;
defparam prom_inst_2.INIT_RAM_02 = 256'hD06BCA20FED06BCAB71AD047C32313D060C2BE1AD056CAB77EDE2A11D12CCAB7;
defparam prom_inst_2.INIT_RAM_03 = 256'h4453C9D074C205C809CD234EE9EBD1F1CD56235E23D03FC32323D060C2B7237E;
defparam prom_inst_2.INIT_RAM_04 = 256'hDAD676CDD21411D09CC2B7D08ECA20FE1A13DE2C11000A0D4E392E38565F534F;
defparam prom_inst_2.INIT_RAM_05 = 256'hC809CD200ED074CD0806D0E9C208E6E17E09000B01D0A3C2FFFEC81BCDE5D0F1;
defparam prom_inst_2.INIT_RAM_06 = 256'h15CD7E6F12C67DD0E6C3C818CDD21F21D0D9CA10E67EC809CD200ED074CD0306;
defparam prom_inst_2.INIT_RAM_07 = 256'hFACA20FE7E23DE2B21C818C3D20021E1C9D0A2D2D6A2CDD1F1CDC815CD7E2BC8;
defparam prom_inst_2.INIT_RAM_08 = 256'hD000C3E1D238CDC818C3D21B21D0D6D6CDEBC818C3DD0021D1F1CDD10EC2B7D0;
defparam prom_inst_2.INIT_RAM_09 = 256'hD47BCDD21611D140D2D471CD2E0EDE2A21D1F1CDC818C3D20B21C000C3D238CD;
defparam prom_inst_2.INIT_RAM_0A = 256'h23D170C24FFE7E23D170C24DFE7E23D471CD2E0EDE2A21D0F1DAD755CDDE2A11;
defparam prom_inst_2.INIT_RAM_0B = 256'h7E2356235EE1D771CDE5DE2A21000401D1A1C3E5200001C00021D170C24EFE7E;
defparam prom_inst_2.INIT_RAM_0C = 256'h15CD79C815CD78C1C809CD2C0EC5C815CD7DC815CD7CE5EB03479A784F934623;
defparam prom_inst_2.INIT_RAM_0D = 256'h0DFE0036D1E3CA18FED1CACA5FFED1CACA08FEC803CDDE2A21D238C3D771CDC8;
defparam prom_inst_2.INIT_RAM_0E = 256'h2BC809CD080EC809CD200EC809CD080ED1AACA2AFE7DD1AAC3C809CD4F2377C8;
defparam prom_inst_2.INIT_RAM_0F = 256'h003A410A0D000A0DC9C818CDD1F821D1C3C323D1AACA0DFED1AACAB77ED1AAC3;
defparam prom_inst_2.INIT_RAM_10 = 256'h44204F4E0D00534B522E002A000D525245000D4B4F00295328454C4946204F4E;
defparam prom_inst_2.INIT_RAM_11 = 256'hFF3EC9F001320C3ED23AC30F3E00D1190049D1200058D0F7004443D08B005249;
defparam prom_inst_2.INIT_RAM_12 = 256'h7AD240CDF579D23ECD000011000021C9F0003A0000D23ECDC9E1C90000F00032;
defparam prom_inst_2.INIT_RAM_13 = 256'h21808011D240CD953ED279CA873E48FEF1D240CD7DD240CD7CD240CD7BD240CD;
defparam prom_inst_2.INIT_RAM_14 = 256'hCDD298C205D23ECD1006D238CDC901D6D282C2B57C2BD079BB924FD248CD4E20;
defparam prom_inst_2.INIT_RAM_15 = 256'h0EC0FEE6D251CD410ED2D3CA01FED254CD480E01AA21C001FED251CD400ED233;
defparam prom_inst_2.INIT_RAM_16 = 256'hFED248CDD248CDD248CDD248CDC9B7F1C818CDD34421F5D2B7CA01FED251CD41;
defparam prom_inst_2.INIT_RAM_17 = 256'h51CD7A0ED2E4CA01FED257CD690E400011000021C0FEE6D251CD770ED2B7C2AA;
defparam prom_inst_2.INIT_RAM_18 = 256'hCD500E020021D248CDD248CDD248CDE1C818CDD34B21E5D324C240E6D248CDD2;
defparam prom_inst_2.INIT_RAM_19 = 256'hCD500E020021DE6232FF3EE1C818CDD35221E5D248CDD248CDD248CDC9B7D254;
defparam prom_inst_2.INIT_RAM_1A = 256'hCD00FF11C5D5000A0D2B32564453000A0D32564453000A0D31564453C9B7D254;
defparam prom_inst_2.INIT_RAM_1B = 256'hD35ACDE5C9002E655C578F2979C93F37001659D373CA00FEDE623AD8E1C1D27F;
defparam prom_inst_2.INIT_RAM_1C = 256'h77D248CD2377D248CD0006C0FEFEE1D27FCDFF0111D246DAD257CD510ED246DA;
defparam prom_inst_2.INIT_RAM_1D = 256'hC1CDAFC954FE7EC041FE237EC046FE237ED93621C9D23ECDD23ECDD397C20523;
defparam prom_inst_2.INIT_RAM_1E = 256'h77897E23778A7E2377837EC946234E2356235EC9130300266C128D0AD3C4CDD3;
defparam prom_inst_2.INIT_RAM_1F = 256'h8F784F8F79578F7A5F877BC947887E234F897E23578A7E235F837EC977887E23;
defparam prom_inst_2.INIT_RAM_20 = 256'h3423C0D41FCDC9F1D3F5CDE1D3D5CDE5D415D2F50FD40BCDD408CDD405CDC947;
defparam prom_inst_2.INIT_RAM_21 = 256'hC9961A2B1BC0961A2B1BC0D438CD232323131313C904C00CC014C01CC93423C0;
defparam prom_inst_2.INIT_RAM_22 = 256'hD458C20D2313771A04D458CAB779000401C967987C6F917DC9B623B623B6237E;
defparam prom_inst_2.INIT_RAM_23 = 256'h13C8B7771AD471C323C837B7C8B97EC9D465C2B1780B2313C0961AC9D458C205;
defparam prom_inst_2.INIT_RAM_24 = 256'hC8CA2AFED4AFCA2EFED4BECAB7D484CD0B0EC9DFE6D07BFED861FE1AD47BC323;
defparam prom_inst_2.INIT_RAM_25 = 256'h203E13D4BEC2D4C4DA04FED4F3CA0BFE79C9D490C20D2313C0BED4A8CA3FFED4;
defparam prom_inst_2.INIT_RAM_26 = 256'hBED4C4CA05203E4702D679D4DBC22EFE1006C8B7D484CD13D490C313D4A6C31B;
defparam prom_inst_2.INIT_RAM_27 = 256'h0D2313C0BE203E1BD4FBC2B71AD4A8C3D490CA2EFE1AC9B7D4DBC20D23D4EACA;
defparam prom_inst_2.INIT_RAM_28 = 256'h7123722373DE1421C8B97E23D518C2BA7E23D518C2BB7EDE1421C9B71AD4F3C2;
defparam prom_inst_2.INIT_RAM_29 = 256'h4B000011C037D293CD00544146000A3631C9F1C818CDD52F21F5D37CC3D90021;
defparam prom_inst_2.INIT_RAM_2A = 256'h2AC818CDD53321C037D3ACCDD8D518CD4FDAC83AEBDAC62AD0D554CDD8D518CD;
defparam prom_inst_2.INIT_RAM_2B = 256'hDE0411D91C01D575C23D19D9103AD90E2AEBD9162AD3BDCDDE0011D91C01D90E;
defparam prom_inst_2.INIT_RAM_2C = 256'h3AD3BDCDDE0811DE0401DE0E22676C8F298F298F298F29DE0C22D9112AD3BDCD;
defparam prom_inst_2.INIT_RAM_2D = 256'hC9AFDD0022005C21DE1222D5C021D526CC36FED93A3ADE1132C33EDE1032D90D;
defparam prom_inst_2.INIT_RAM_2E = 256'h7B56235E19D90011290026DE1D2AD5ECDAD506CDD3E5CDDE0021D3CDCDDE1E21;
defparam prom_inst_2.INIT_RAM_2F = 256'h1D21D637C2B7DE183AE5C9DE1F22DE1D22676FAFC9DE1D22EBD5ECCA3CA207F6;
defparam prom_inst_2.INIT_RAM_30 = 256'h57987E235F917EDE1D21000201D44FCDDE1921DE0811C937E1D60AC2D440CDDE;
defparam prom_inst_2.INIT_RAM_31 = 256'h235EDE1921DE18323DDE103AD5C0CDD402CDDE1921DE103A47987E234F987E23;
defparam prom_inst_2.INIT_RAM_32 = 256'h6FAFD8D64ACDDB0021D65FC2B7DE253AD37CC3D5F6CDC9E1D41ACD2B2B4E2356;
defparam prom_inst_2.INIT_RAM_33 = 256'hECCDD690C2B7DD013AD5C919DB00112929292929DE2532AFD669DA10FE3C0026;
defparam prom_inst_2.INIT_RAM_34 = 256'h2532AFDE1832AFD44FCDDE1D21DE2611D69AC3DE0E3AD44FCDDE1921DE0411D5;
defparam prom_inst_2.INIT_RAM_35 = 256'h8ECDE5D5D6A2CAE5FE7EC837B7E1D6ACC20D23B6AF200EE5D8D1D650CDD5D1DE;
defparam prom_inst_2.INIT_RAM_36 = 256'h13DD0132D6E3C25CD61AC956235E1900051146234E19001411D6A2C3C8D1E1D4;
defparam prom_inst_2.INIT_RAM_37 = 256'h0B11E5D709DAC1D676CDD5E5D1EB13121BD6E4C25CD613D6F2CAB71AD5C8B71A;
defparam prom_inst_2.INIT_RAM_38 = 256'h237EDD0021D170237123722373DE2621D6C7CDC5D5D8D13F07070707E17E1900;
defparam prom_inst_2.INIT_RAM_39 = 256'hC3DD0032D733C25CFE00367E2BD74EC22EFE1A13D742C22EFE1AD71FC2B77E47;
defparam prom_inst_2.INIT_RAM_3A = 256'hCDD8D676CDDE2322000021C9D6E3C2B71AD1D47BCD235C36D74BCA5CFE78D74E;
defparam prom_inst_2.INIT_RAM_3B = 256'hD448CDD798CAB57CDE232AE5C8B178C9DE1832AF70237123722373DE1D21D6C7;
defparam prom_inst_2.INIT_RAM_3C = 256'h21C5D7B4D202FE78E5C1D452CDEBDE212AE5D448CDE14D44DE232AC5D1D7C6D2;
defparam prom_inst_2.INIT_RAM_3D = 256'hC1D64ACDC5E1DE2322000021C9D771D2E1C1D64ACDDE2122DB0021DE23220200;
defparam prom_inst_2.INIT_RAM_3E = 256'h000000000000000000C9EBDE2122EBD452CDE1EBDE212ADE2322D771C30505D8;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ad[12]),
  .CLK(clk),
  .CE(ce)
);
MUX2 mux_inst_2 (
  .O(dout[0]),
  .I0(prom_inst_0_dout[0]),
  .I1(prom_inst_2_dout[0]),
  .S0(dff_q_0)
);
MUX2 mux_inst_5 (
  .O(dout[1]),
  .I0(prom_inst_0_dout[1]),
  .I1(prom_inst_2_dout[1]),
  .S0(dff_q_0)
);
MUX2 mux_inst_8 (
  .O(dout[2]),
  .I0(prom_inst_0_dout[2]),
  .I1(prom_inst_2_dout[2]),
  .S0(dff_q_0)
);
MUX2 mux_inst_11 (
  .O(dout[3]),
  .I0(prom_inst_0_dout[3]),
  .I1(prom_inst_2_dout[3]),
  .S0(dff_q_0)
);
MUX2 mux_inst_14 (
  .O(dout[4]),
  .I0(prom_inst_1_dout[4]),
  .I1(prom_inst_2_dout[4]),
  .S0(dff_q_0)
);
MUX2 mux_inst_17 (
  .O(dout[5]),
  .I0(prom_inst_1_dout[5]),
  .I1(prom_inst_2_dout[5]),
  .S0(dff_q_0)
);
MUX2 mux_inst_20 (
  .O(dout[6]),
  .I0(prom_inst_1_dout[6]),
  .I1(prom_inst_2_dout[6]),
  .S0(dff_q_0)
);
MUX2 mux_inst_23 (
  .O(dout[7]),
  .I0(prom_inst_1_dout[7]),
  .I1(prom_inst_2_dout[7]),
  .S0(dff_q_0)
);
endmodule //t20k_rom
