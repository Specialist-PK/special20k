//Copyright (C)2014-2024 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.10.03 (64-bit)
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Mon Dec  9 18:59:07 2024

module t20k_romram (dout, clk, oce, ce, reset, wre, ad, din);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [12:0] ad;
input [7:0] din;

wire [29:0] sp_inst_0_dout_w;
wire [29:0] sp_inst_1_dout_w;
wire [29:0] sp_inst_2_dout_w;
wire [29:0] sp_inst_3_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

SP sp_inst_0 (
    .DO({sp_inst_0_dout_w[29:0],dout[1:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1:0]})
);

defparam sp_inst_0.READ_MODE = 1'b0;
defparam sp_inst_0.WRITE_MODE = 2'b00;
defparam sp_inst_0.BIT_WIDTH = 2;
defparam sp_inst_0.BLK_SEL = 3'b000;
defparam sp_inst_0.RESET_MODE = "SYNC";
defparam sp_inst_0.INIT_RAM_00 = 256'hE552E0B2CBC8D6F83577E2D9F6E2A8C82655557A2935555C7A07A41500FEAF4F;
defparam sp_inst_0.INIT_RAM_01 = 256'h9A27A9E6589E2499EA78B21F2041252C2CBA09959B4EFAD55095DDCDD9C88A74;
defparam sp_inst_0.INIT_RAM_02 = 256'hA77EED9518E7B6CBC8104017E96657E966597F96A1727C957E966497F9EA177B;
defparam sp_inst_0.INIT_RAM_03 = 256'hD7CB2696F9AADA15E6E2E9EECA9BAB685AF2B795FE551D89BD4595495546977E;
defparam sp_inst_0.INIT_RAM_04 = 256'hE5169BBB687B62F97E67EA5D1C958B4BFDBB1860A5EF65EA66EEDA1E6A4EEE3E;
defparam sp_inst_0.INIT_RAM_05 = 256'hBE7EF246FB2E991E8A157AE1B5BD0FC955564FA55CBF287B2FC8FBD5647D5D96;
defparam sp_inst_0.INIT_RAM_06 = 256'hB6C940004A225209FC13A3CBE5F94789561563763EBDF8A3476ACB22CBE172AC;
defparam sp_inst_0.INIT_RAM_07 = 256'hBF780157A41F9B07FA9BE2D54FF957EE96FBBA6CFEFAA7AEDB6D77ED8A2DBF9D;
defparam sp_inst_0.INIT_RAM_08 = 256'h0020021DB7EF8EA09BD7ED4117D04D0F342E4637E9D20BE42CDFD2FD2FD2FBF4;
defparam sp_inst_0.INIT_RAM_09 = 256'h00CEE4E40044E4E70089F9DE0088387600F0817900600D91316F83000CFA0C1A;
defparam sp_inst_0.INIT_RAM_0A = 256'h0024000000C0000000C0019002A02002002A19283C24098C2BBA002A00000000;
defparam sp_inst_0.INIT_RAM_0B = 256'h00960260033020020000000009D625960027258325632BAA25A7309620002576;
defparam sp_inst_0.INIT_RAM_0C = 256'h25561755155D340018092555200215D537060083308325562406259617582376;
defparam sp_inst_0.INIT_RAM_0D = 256'hC00000182AAA0600200230A70025162525550295255500032586189619560096;
defparam sp_inst_0.INIT_RAM_0E = 256'h255615D5155D15571C0D1575157516250007035C32A31EAA1EAA258317562556;
defparam sp_inst_0.INIT_RAM_0F = 256'hFFFF15D51D5525D6355525961555258025961595009520072406009615D71557;
defparam sp_inst_0.INIT_RAM_10 = 256'hA9EE288E22B86259AE217D565E4B37EB7607D2CB0477D30638E79E3EF38FFFCB;
defparam sp_inst_0.INIT_RAM_11 = 256'h76441F9107644A5752E717E7E415FEFE50547E50BA38BB6E2A92E698AA188AE4;
defparam sp_inst_0.INIT_RAM_12 = 256'h9F6FB6F41F9765FBD9AF4B757114799579076EBED5B9AF779657655465117B90;
defparam sp_inst_0.INIT_RAM_13 = 256'h6971979071C5E5E6F4A9E6F7BECB9C75975F9AD8FA8B5F90556BFAAD2D145907;
defparam sp_inst_0.INIT_RAM_14 = 256'h72526F5971AC1CA5D41FA5E41EA5C7D88D1E85FBCBEBF4BF4B5BFEADE6B5C6AF;
defparam sp_inst_0.INIT_RAM_15 = 256'hAFC8DC6C6C7C4C55C6B9E79AFC6AEC6A716EC6B9EA2D4B9B6B1E71C65D7E4155;
defparam sp_inst_0.INIT_RAM_16 = 256'h656D9726CF8A2C55F361287A127C97A0CF61DF6C8DDBE6C8BD472712EAF1317E;
defparam sp_inst_0.INIT_RAM_17 = 256'hF7A65ED0F6171E9C1CB6F07A7D957E77ACE6E9BCB69435EB97A557F1F9147E57;
defparam sp_inst_0.INIT_RAM_18 = 256'h14559656512FC35F65965965814EA3FC368BC352F0D7D965604A659656DF7755;
defparam sp_inst_0.INIT_RAM_19 = 256'hF87647E47647CAC47F652B43658686E389D0BDA2055DF18D0C1E138D76050597;
defparam sp_inst_0.INIT_RAM_1A = 256'h520E1F499E2000000079BDC51715227A2E89B92A889DFF555D58868172DBF876;
defparam sp_inst_0.INIT_RAM_1B = 256'h8BA26E9AA62519F7FF67D5753D3F55625AA9F659607DF5574E1287A12D236749;
defparam sp_inst_0.INIT_RAM_1C = 256'hFB8B8BAABB2A5561652CEF4E86FF658B43659620584A7E10BA7975498749E61D;
defparam sp_inst_0.INIT_RAM_1D = 256'hB6EABAA53642C9656529798890E54BA6AE787E1FFD5878695639BBB685B93BB9;
defparam sp_inst_0.INIT_RAM_1E = 256'h8000011157160E2F0CB1B4A179F18696165A29572076727F2EBE7FBF88890552;
defparam sp_inst_0.INIT_RAM_1F = 256'h04C7050121041441C618500024FC6079F9136109A6F84D849819A089A0C49854;
defparam sp_inst_0.INIT_RAM_20 = 256'h34245E756ECFF0BE388EE3FC2A2BA94BAD41745A05105D19CA927421F2C51049;
defparam sp_inst_0.INIT_RAM_21 = 256'hA2BB43854AA5516C5BA4B06D18A1481E14812189934EE351A9842CA2B84998BF;
defparam sp_inst_0.INIT_RAM_22 = 256'hBB9D5A415D0414AAD2EB49AC5AA46D69369485AA550ED0E10D843B4A70D155AC;
defparam sp_inst_0.INIT_RAM_23 = 256'h26494145FDA66B9BC52148526A96C5FC62789AE688DA63D4545114915147F8FB;
defparam sp_inst_0.INIT_RAM_24 = 256'h4185A6E2616121E1A15A410508295402E462AF8514030CC90E4FA21A47C7118E;
defparam sp_inst_0.INIT_RAM_25 = 256'h5A89AD60412A5EBAA186185D0716E6958A95AE684991A52B62692856A931EE18;
defparam sp_inst_0.INIT_RAM_26 = 256'hE5493D5F27E2A85B4D527A3268C963784A1AB907961861784A18618507D72286;
defparam sp_inst_0.INIT_RAM_27 = 256'hCF7EFDCBDBEBF9CBDBEBF9BBB9F226C75D286E2B9969A7E7E1F848A6DD6AB5AA;
defparam sp_inst_0.INIT_RAM_28 = 256'hCF87CF19193F290909FE02D05C356EEE6BCAF01FFF40004C30D5D5D519CD0457;
defparam sp_inst_0.INIT_RAM_29 = 256'h7C8B3B830AA739CA824BA4EA23070F2F2CA088EE509F20B82A3A8AC1E78E1A3F;
defparam sp_inst_0.INIT_RAM_2A = 256'h85159526B6B585168174F111E2EA1111C13B418A54175CD17BE11B4AB4BA178E;
defparam sp_inst_0.INIT_RAM_2B = 256'h5BB896E9BF66D22EEE514A6499D61D697481A91629A9BA25B5861AB3777625B5;
defparam sp_inst_0.INIT_RAM_2C = 256'h18B595C5559B9882F29C6EE6CD9527EEE96262449962CBCBCBDA524D96176A06;
defparam sp_inst_0.INIT_RAM_2D = 256'hD766957EE22EAE4ED6B8A6E45B906B1495A9A3D89EC918566E2CD969AEA36585;
defparam sp_inst_0.INIT_RAM_2E = 256'h0724B9118B37BE5B4A6E05BB9372F88ED2F88AFAABEAAFBBE4537BE9B547FF64;
defparam sp_inst_0.INIT_RAM_2F = 256'h000000000000000000001E6C979AEDD4695B81765A66C6E85CA852799054B97A;
defparam sp_inst_0.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_1 (
    .DO({sp_inst_1_dout_w[29:0],dout[3:2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:2]})
);

defparam sp_inst_1.READ_MODE = 1'b0;
defparam sp_inst_1.WRITE_MODE = 2'b00;
defparam sp_inst_1.BIT_WIDTH = 2;
defparam sp_inst_1.BLK_SEL = 3'b000;
defparam sp_inst_1.RESET_MODE = "SYNC";
defparam sp_inst_1.INIT_RAM_00 = 256'h8EA1E27847F7C7C72AB761E2BC103FF8639560B600A555503A03480505303F00;
defparam sp_inst_1.INIT_RAM_01 = 256'hCAF1ACAB3AC6B2BC2B18FE03C2030F231F3911F8E78C7AE0031D439438EA4444;
defparam sp_inst_1.INIT_RAM_02 = 256'hB3F0BC952C2BFACCF080C00CE4C7CCE4E3F4C44A3CC1103CCE407C4C440FCC1B;
defparam sp_inst_1.INIT_RAM_03 = 256'hC4D3E2123401C87104F1C8CFC8B28721C2760F540F603C0D100D5A01600113F0;
defparam sp_inst_1.INIT_RAM_04 = 256'h8C3523C721FC23F9B03B03103D20D745561BFC811E5F210044F1C87D8ABBF48D;
defparam sp_inst_1.INIT_RAM_05 = 256'h86BE7663F3020C338C30F8C30C7802FA55801FA58F2BE3FFC0F9B78603786FA0;
defparam sp_inst_1.INIT_RAM_06 = 256'h724D40008C83218C2002C0CBC8030F4E00B5482C8E3C13C80C2BD3C1F80202BF;
defparam sp_inst_1.INIT_RAM_07 = 256'hF1FC02004DBC0E6FC3456B5501FA0B2019C3C0B330C078C6C722F0685A3CB76C;
defparam sp_inst_1.INIT_RAM_08 = 256'h020800EC88FF1EB8BC7B22DB7FC510601E3F9C5C0EB2D4F941747B47BC7BC11E;
defparam sp_inst_1.INIT_RAM_09 = 256'h00FA550000CA550200AB9D9200F5F01900FC26CC00E88AAC330703E0033E0C06;
defparam sp_inst_1.INIT_RAM_0A = 256'h02403C0000C027C005D405D4240606A4004531E9024A1DDD2BBA002A11550000;
defparam sp_inst_1.INIT_RAM_0B = 256'h110324060330062427CF3C3C30C330C32A4330C93033032430433243355D3243;
defparam sp_inst_1.INIT_RAM_0C = 256'h300300600058300001903000355700C0300300C330C33AAB300330C303093143;
defparam sp_inst_1.INIT_RAM_0D = 256'hC0000009300300603AAB32C315600260254016803000155730C301C3310300C3;
defparam sp_inst_1.INIT_RAM_0E = 256'h340700C000582AA901900241024002600003175D30C30EA90C0030C3030305D4;
defparam sp_inst_1.INIT_RAM_0F = 256'hFFFF00C00D55304335543043258030C030C305D409803557300300C309C30003;
defparam sp_inst_1.INIT_RAM_10 = 256'h8EA79AFA7EAFEFDBFE7CF3EFFC24AF8F3083C82C0B8A200ACF3CF3CA00E04124;
defparam sp_inst_1.INIT_RAM_11 = 256'hF6AFFDABFFEAECC8D7D34BAB8BF81EFBBFE6C378FF48BE23C9E678AF6FAAF638;
defparam sp_inst_1.INIT_RAM_12 = 256'h87ADB4080C0701F2F230A49C22BAC6BB38238DF4989AC6A0FFB6BF8AFFAB6E6F;
defparam sp_inst_1.INIT_RAM_13 = 256'h2FF0FFC5F0C28E8B1ECE8B1FF0C6BC30FF0F2A7A3CA98C23B568F2A792BAEB23;
defparam sp_inst_1.INIT_RAM_14 = 256'hBE8DDC1FFC83FFBFE3FCBFD3FEBFC33B172EBBCAF2E11EF1ECBA02A68AF0C2A7;
defparam sp_inst_1.INIT_RAM_15 = 256'h808970F0E0E0F0F00DEFBEF900E27C28C3B30DEFF22606B0FF0AF0C3FC308ED5;
defparam sp_inst_1.INIT_RAM_16 = 256'hA03E2E8F3B3F3C166C3BBEFFBB6BAE8BB03BD76B97D2EF8AC7DA0C33F803C3F2;
defparam sp_inst_1.INIT_RAM_17 = 256'hCE4F7FF07ABF4B13F57AAFECEE956043C34BF9DC3AFE5CF38788003CE3EDF656;
defparam sp_inst_1.INIT_RAM_18 = 256'h07B8EFFFFDD025CCFFFE4EFFFF72EE025CF025CD09733FFF7FFAB8EFF7B02C00;
defparam sp_inst_1.INIT_RAM_19 = 256'hD0B4CF0CF0CCC2C3CCFFC065FBEFFAFD8ECF9DB1FE220E17F3378E977302FCFF;
defparam sp_inst_1.INIT_RAM_1A = 256'hF4B3BDCBF6B0000000C8C7C17706119747D8F76BD8E3036ABBEBEF80B2CAC9F6;
defparam sp_inst_1.INIT_RAM_1B = 256'hD1F63DEAFA383B1D55EC77878B81CFEBEAF71FBFFFF3EE01D3BBEFFBBB65F8D2;
defparam sp_inst_1.INIT_RAM_1C = 256'h3D2BC72C3F22D6077790F1CFFFCCFFD065FBFF1FEECFC3B8FF8FF884EF4653BD;
defparam sp_inst_1.INIT_RAM_1D = 256'hFECAF2BA1F1BFA3737BDFDC8C3798576BDBFE7FFFE0EEEEFD4813C721EDAEF7D;
defparam sp_inst_1.INIT_RAM_1E = 256'hC0000330F403BC7E0C36FCA022B2EEE3BB6B2E03C23C70C13EBCC181AC48015B;
defparam sp_inst_1.INIT_RAM_1F = 256'h0C0C0EEB23CE34D30C34C00035D48022BB30440AF7E8C110AECCE0B860C38438;
defparam sp_inst_1.INIT_RAM_20 = 256'h4846B3A0D30C001328CA61000E19F839CC481EBFAF0AC833078B5CC281420ACC;
defparam sp_inst_1.INIT_RAM_21 = 256'hA3CE2800804C39FA7F1C4ACC287ACC71ACC79224E200FAD09710C4E38F0BEE73;
defparam sp_inst_1.INIT_RAM_22 = 256'hC4C4DE040100003F00FC03F13FE025F86C4013FE03A0800B002E8205EA300CC4;
defparam sp_inst_1.INIT_RAM_23 = 256'h22CBAB2000AF29C8ABBACEBB2AF22BC6F10ACAF2AE3E084E7A78AFD9F9F61AC4;
defparam sp_inst_1.INIT_RAM_24 = 256'h000DCA7B03C3C3838363C002080F8800F80F23C2202110824FC232304EC89E4F;
defparam sp_inst_1.INIT_RAM_25 = 256'h3B18C7B000343712CB2CB2E4AC44630CCD0CC231EC80C330C84F12E101E28CBC;
defparam sp_inst_1.INIT_RAM_26 = 256'h2D8DDEAD1823CA03CC52E142C50B1491CC0C3CAC04B2CB91CC02CB2CAC84412C;
defparam sp_inst_1.INIT_RAM_27 = 256'hEF9EDA6CEC6CCE6C6C6C4E4C4E01CE1C3E7C331CE48F3C444B12C4F0FC061CC6;
defparam sp_inst_1.INIT_RAM_28 = 256'h259025AE50A01A6163065A6126F391139A86A1B00093139041F81C1D51DB6D79;
defparam sp_inst_1.INIT_RAM_29 = 256'hC0CE61984BE9631AD64D198F195C405231C59D2BA43036BDAB7BDE57BB4B8E60;
defparam sp_inst_1.INIT_RAM_2A = 256'hD2C53A2BA98FC2CBAB404F9BEAA6179B8010C44922B713200034AC62C62F4990;
defparam sp_inst_1.INIT_RAM_2B = 256'hC51E9BCF1FBC9EC593A087E7971F03FCBC0CC105DEAC0F0B8FE34F1FBBBBC88F;
defparam sp_inst_1.INIT_RAM_2C = 256'hF41C9A82AAD368F1F9B81C7631786EB13E38F24D3E326CEC6CCFC01FE389184F;
defparam sp_inst_1.INIT_RAM_2D = 256'h85A1752094D126663043693844E11081F549F94731CD84D34F8DFF3463E7F8D1;
defparam sp_inst_1.INIT_RAM_2E = 256'h6DA7C98AE30003C5E5F0024186CD6BE73043C79CF843E71D3C0000345D635538;
defparam sp_inst_1.INIT_RAM_2F = 256'h000000000000000000002B0932CB04161B4C009006F08300150E44EC96CDC914;
defparam sp_inst_1.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_2 (
    .DO({sp_inst_2_dout_w[29:0],dout[5:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5:4]})
);

defparam sp_inst_2.READ_MODE = 1'b0;
defparam sp_inst_2.WRITE_MODE = 2'b00;
defparam sp_inst_2.BIT_WIDTH = 2;
defparam sp_inst_2.BLK_SEL = 3'b000;
defparam sp_inst_2.RESET_MODE = "SYNC";
defparam sp_inst_2.INIT_RAM_00 = 256'hCEB2900E903B130B2AA0A92F8F037F385BF188CE23CAAAA00E0CEC2200333FC0;
defparam sp_inst_2.INIT_RAM_01 = 256'hC4301CC720C0720C4302CE00E084080323E007F3CAC8CF09300AC8EC8D380C18;
defparam sp_inst_2.INIT_RAM_02 = 256'h303333A3088FCB0438210004805FC48457F8484D3C4210204809FC84805FC411;
defparam sp_inst_2.INIT_RAM_03 = 256'h8C3CB00030C2CC4300FFCCCFCC400B3108CF03088788C3CE001100100C832033;
defparam sp_inst_2.INIT_RAM_04 = 256'h804423CF3130032C33733330C3C8CAE00334300820EB33040CF3CC4C818CE80E;
defparam sp_inst_2.INIT_RAM_05 = 256'hC886CFDB2CF04CC00CC30B8800CA123BC62C50BE03A8E310EA3BBCA084CAA280;
defparam sp_inst_2.INIT_RAM_06 = 256'hB34100001813C94F2020CC3CB00013101809002003BE10C020CF3CB02C80C8F2;
defparam sp_inst_2.INIT_RAM_07 = 256'hE33C001C400CCB01CCC93074103C18F0113FC0730F8CBCFF4B300C0C853CC3B4;
defparam sp_inst_2.INIT_RAM_08 = 256'h018000E28CF3C8300CC8A30C20414E32303308208CF3C4F0488CC34C34C32A30;
defparam sp_inst_2.INIT_RAM_09 = 256'h0040000000BFFFFF00EFEABA00BEAFBE00EABEBF00042450381059E0000F2687;
defparam sp_inst_2.INIT_RAM_0A = 256'h0400000000400000004001100000000000000500040504100110000000000000;
defparam sp_inst_2.INIT_RAM_0B = 256'h0004000001100040000000001014051400010550041501400401140400000554;
defparam sp_inst_2.INIT_RAM_0C = 256'h0554155515551555155505000000155505541555155510010554155515500554;
defparam sp_inst_2.INIT_RAM_0D = 256'h4000001000000004000014010005140505550015055500010414155505541555;
defparam sp_inst_2.INIT_RAM_0E = 256'h0554155515551000155515551555140515550154155514000555155515541555;
defparam sp_inst_2.INIT_RAM_0F = 256'hFFFF005505550404155504041555155515551515101500050554155510141555;
defparam sp_inst_2.INIT_RAM_10 = 256'h1C4711CC730C8320C8320000418C00AF8A0BF10000010400C10410410400C30C;
defparam sp_inst_2.INIT_RAM_11 = 256'h0A108184206104000014A0A0A0865B6C82188880CC400C8730C8330C4330C031;
defparam sp_inst_2.INIT_RAM_12 = 256'h6C718AAC22ACA81A18768C12EC410C4105387FC6A13C8F22108204C104C42202;
defparam sp_inst_2.INIT_RAM_13 = 256'h310E10210138400730C00733CF8C41421023CCF10F13C1A801843C4F30410434;
defparam sp_inst_2.INIT_RAM_14 = 256'h0E233CA10E30808428828418808428020850802A0A0A30E30CC0184C0D01384C;
defparam sp_inst_2.INIT_RAM_15 = 256'h320081313131313912C000002104F38C047012C03CCF0E123CE101384086A006;
defparam sp_inst_2.INIT_RAM_16 = 256'h4830F083822F0288C400003000213C0F12000C71081C4300CC004043C304C4C6;
defparam sp_inst_2.INIT_RAM_17 = 256'h00C484700320E1080003A200E0F18C28280F0A01C3002208283E4EC20F200218;
defparam sp_inst_2.INIT_RAM_18 = 256'hA000204C4C00820000100204C808C30820CC8231208000043208F02043128493;
defparam sp_inst_2.INIT_RAM_19 = 256'h0A82102102100C2080003202080201F06F2330C420C8F2080080F208C3002210;
defparam sp_inst_2.INIT_RAM_1A = 256'hC4F80320C03000000026CC0054A8D7345314D81F16C0422A8822C302030A0802;
defparam sp_inst_2.INIT_RAM_1B = 256'h14C53607C5B0C8300020C040888B100301C43081320030931000030008420413;
defparam sp_inst_2.INIT_RAM_1C = 256'h3A03FF303F3108C4C8307307108000320208134200204800CC41023700DCDC03;
defparam sp_inst_2.INIT_RAM_1D = 256'hCF01C03C30DF3CC808023026CC3F3001321334C00440000204033CF3120633A0;
defparam sp_inst_2.INIT_RAM_1E = 256'hAAAAA83AAFBAEBEA2EEEAA82AAE8000004040F90E380081B43C01B5B73114867;
defparam sp_inst_2.INIT_RAM_1F = 256'h0D4C4E08830C30C30C30C2AAAABEBEAAE03BBAABBAA0EEEABBAE82EA82EAAAE8;
defparam sp_inst_2.INIT_RAM_20 = 256'h11C008A7199CA63B62D8D4258D53D963D696600C11211E508DAC710F2301211E;
defparam sp_inst_2.INIT_RAM_21 = 256'hCBE6844A1961C1384E4D811651B021C0021C060AC018F1275C554D0B56403B54;
defparam sp_inst_2.INIT_RAM_22 = 256'hE66726806280270F9C3E70F9C869D51971545C869C11201C427045952112710D;
defparam sp_inst_2.INIT_RAM_23 = 256'h30000479098363D88000200062F6002C3361D0740C069C704C4C0201313A0712;
defparam sp_inst_2.INIT_RAM_24 = 256'h8141DC33D0D0D0D0D0F70108CC1C2033F33370C5061701042004620500098020;
defparam sp_inst_2.INIT_RAM_25 = 256'h4C60D48042394C72D041040F112DC3500E50143500A0D407141C470143E7D102;
defparam sp_inst_2.INIT_RAM_26 = 256'h520A52CF15C36D870D102D103440D1351026FE11690410351024104211298241;
defparam sp_inst_2.INIT_RAM_27 = 256'h30D34C0E0E4E4CCECECECC2264429041087C3B0EDE1C7142D0B400F9CC515111;
defparam sp_inst_2.INIT_RAM_28 = 256'h4F5C8F3C63C91450509D14F009E73BBB164591CA95001138E143725257104100;
defparam sp_inst_2.INIT_RAM_29 = 256'h24ED735852D35098D02C1D4B43415161B5C44DC3C509363D0B62DCD0019F6D72;
defparam sp_inst_2.INIT_RAM_2A = 256'h45473574A59C45448478D8541392545401350403CC46B712EED63E53E53D635C;
defparam sp_inst_2.INIT_RAM_2B = 256'h6735E165AA1698E3D951896650612416248659263DF5CD74DC4504A88889259C;
defparam sp_inst_2.INIT_RAM_2C = 256'h8534D146AA6E65F2A50494DB71C252899597D74105971E1E5E5D601059139041;
defparam sp_inst_2.INIT_RAM_2D = 256'h1911C6655855CD4D53615194121158190962F3E60BA25515B979059951341645;
defparam sp_inst_2.INIT_RAM_2E = 256'h414F6A3C5EEEED64171A0863572741F41371CF90B542D53CB49EEEDA405700B4;
defparam sp_inst_2.INIT_RAM_2F = 256'h0000000000000000000009A94A69A7011026821D841A49A0874F8526A4206851;
defparam sp_inst_2.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_3 (
    .DO({sp_inst_3_dout_w[29:0],dout[7:6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:6]})
);

defparam sp_inst_3.READ_MODE = 1'b0;
defparam sp_inst_3.WRITE_MODE = 2'b00;
defparam sp_inst_3.BIT_WIDTH = 2;
defparam sp_inst_3.BLK_SEL = 3'b000;
defparam sp_inst_3.RESET_MODE = "SYNC";
defparam sp_inst_3.INIT_RAM_00 = 256'h7010402C6C3D604D301AC3B1EC3EEDB3F37FFFECCE4FFFF02CC2C00F0DF08733;
defparam sp_inst_3.INIT_RAM_01 = 256'hF73DCF33CCF33CCF33CCECDEC03333DD0B13FFDE787BAC7FFEC0774777B0370F;
defparam sp_inst_3.INIT_RAM_02 = 256'h0EF00B3F3BB5EC7BB00CC0374F7F774F736374F33770DCCF74F3F4374F3B77DC;
defparam sp_inst_3.INIT_RAM_03 = 256'h7BB2CFCFF3F3C37EF3FFC3FFC37DCF0DFFACEF3FB4FF7B13EFEC3FEC7FCDCEF0;
defparam sp_inst_3.INIT_RAM_04 = 256'h73B0DFCF0DF37BB3F08F08EF7B3F71AC01CC30F7CFF30EF333F3C37C730CC73C;
defparam sp_inst_3.INIT_RAM_05 = 256'h37ECACF3B2CCEF7DEFBEECB7EC2CDFB1FFFFB2CFFB02CED2C0B032CFFB2CFB3F;
defparam sp_inst_3.INIT_RAM_06 = 256'hF043C000CFF7F3DFCC0EFFB2CFDCEF03FFFFFFEFFB3CDEFFEF33B2CBB333F73B;
defparam sp_inst_3.INIT_RAM_07 = 256'h1DF003FFF3BC0DEDC0CD107FEDB3FACEC0B33B3EECBBF7B94F0FDBB8F7BC11D4;
defparam sp_inst_3.INIT_RAM_08 = 256'h00BF33FB37CB373CCF3ECFF3CECE34CCCF35F3CC079E73CF333770770770B1DC;
defparam sp_inst_3.INIT_RAM_09 = 256'h002A00000000000000155555001555550041555500020002015550000FEC0438;
defparam sp_inst_3.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_10 = 256'hDFB7FDF37DDFB7EDF37FF7DF3D33DE872CC1CFFF0FBEFB0F7DF3EF7CFFFF7CF3;
defparam sp_inst_3.INIT_RAM_11 = 256'hE8CF7A33DE8CFF3CF0F28E8E8F7311473DCFB3FCD73EDF77CDF37EDF37EDF77E;
defparam sp_inst_3.INIT_RAM_12 = 256'h868A28000A3E8FA3A310F3DF477DF37D28028C68FDE739FCCF3FFB7CFB73C47D;
defparam sp_inst_3.INIT_RAM_13 = 256'hCCE8CF8CECA3F3FFDC03FFDF2C833B2CCF8B3B9FECFE7A17BFF3B339CF7DF702;
defparam sp_inst_3.INIT_RAM_14 = 256'hECF00C3CF8DF7A33E37B33E37A33D37DF35A3BB3A3A1DC1DC3FCC33BF86CA33A;
defparam sp_inst_3.INIT_RAM_15 = 256'hFCCF3FDFDFDFDFDFFF33CF3FCFFF9A3B3FC0FF33B3B9C0EC368CECA33E285EFF;
defparam sp_inst_3.INIT_RAM_16 = 256'hBF3A13730DCD093F73FF0FD3F0CCE779CCFF768CF3A373DCF35F33F0CDFF7F68;
defparam sp_inst_3.INIT_RAM_17 = 256'hDFF3F44A68EF4FC334E80DFF0A3FFB0E8339A35A28DFCFA28E87F468A1FD68FF;
defparam sp_inst_3.INIT_RAM_18 = 256'h4FBFCFB7B7DC3CFDF7ECFCFB77F78CC3CC733CDCCF3F7DFBDDF39FCFBDECFBFF;
defparam sp_inst_3.INIT_RAM_19 = 256'hA168CE8CE8CCA093BDF7EC3CF3FC3F7FCD6EEA10DFF30EF3EFB67EF3D903DFCF;
defparam sp_inst_3.INIT_RAM_1A = 256'h7793F5ECFB30000000DCF3A35E4F33CF37CDDF73CCF3318033CCF300E8A3A168;
defparam sp_inst_3.INIT_RAM_1B = 256'hCDF377CCF73FBFCD00FF3FFFB3B1FFF3FCF7CF3EDDF7CFFDDFF0FD3F037CF7DE;
defparam sp_inst_3.INIT_RAM_1C = 256'hF1DFFF0EFF0DFFF7F7CF3CF3DF3DF7CC3CF3ED0DFFC333FCD77CF4CFFDCF3FF7;
defparam sp_inst_3.INIT_RAM_1D = 256'hECCCF337CFFFB3FFFF0FD3FCF737CCFF33DED7B007FFDFDEFF7CFCF0DDEC331E;
defparam sp_inst_3.INIT_RAM_1E = 256'h0000000155155555005554005553FC3FF0F0CDFEC33333010B330101102083FE;
defparam sp_inst_3.INIT_RAM_1F = 256'h0141405100410410410410000554545550015505555005545555401540055454;
defparam sp_inst_3.INIT_RAM_20 = 256'h5F7331FFD1330DE1DCF78DC378DE70CE70F0EF30CF0CFCCC0300CF3900030CF4;
defparam sp_inst_3.INIT_RAM_21 = 256'hF34C33C3FBEFFCD33537FCF0FCDCC370CC370FCF403BFCFFF7C3BBB30C004055;
defparam sp_inst_3.INIT_RAM_22 = 256'h447DFC00EF030DDD3774DDD370C3FDF0DF0DF70C3FCF0CF3CFCF3C3FFCF0FF3B;
defparam sp_inst_3.INIT_RAM_23 = 256'h0400F3F3F3B3EE7B330CC330ECDEF34730FCFF7FCF3C33DF3737CC3CDCDF1964;
defparam sp_inst_3.INIT_RAM_24 = 256'h28DE3787F777777777DCC003C033FC30CF00CC0C1C1F17854505400541411545;
defparam sp_inst_3.INIT_RAM_25 = 256'h74FCF74400FF74EEF7DF7DFBCF4FB3DD3FDD3F3DD08CF74CFB330CF3EE4DA774;
defparam sp_inst_3.INIT_RAM_26 = 256'hDFC158700773D3FDCCF00150054015EDD00D33CF4F7DF7EDD00DF7DFCF4F37DF;
defparam sp_inst_3.INIT_RAM_27 = 256'h965967646464676464646744470048FFFB7771DC70F3CFB0771DC3FF7C37DD37;
defparam sp_inst_3.INIT_RAM_28 = 256'h393732E7DE40E3DCDC0437903659E221E0380F3000CCCCC30F3FFFFFCF33CF3D;
defparam sp_inst_3.INIT_RAM_29 = 256'h0380FE3BECCEFC3FBF0137F30EECECEC03BFCFF37EC0EECFF3ECFBBB0FF7DCDC;
defparam sp_inst_3.INIT_RAM_2A = 256'hC30DC30C3C3BC30C33C33BF37CFCF7F340CEC5403F3C3DF04470E4CE4CE70E3F;
defparam sp_inst_3.INIT_RAM_2B = 256'h0CEC3F0C16F0FF235130030FF3FF0FF0EC04C3CCCF0C330C3BC30C1622230C3B;
defparam sp_inst_3.INIT_RAM_2C = 256'hFEEC3CC000C2DCC06F7C37B0DFFFCC111C3030FF3C30646464670037C30CF3DF;
defparam sp_inst_3.INIT_RAM_2D = 256'h0F3F7FF03F73F8F830FDCD1004403BFFBFEFDCBEC283FDFF0B0B7C30EF0DF0C3;
defparam sp_inst_3.INIT_RAM_2E = 256'hDFB9C3E7C244470FFDF003FE3DC4DDDDF0CDC13730DCCCE51C344470FFFC00D0;
defparam sp_inst_3.INIT_RAM_2F = 256'h000000000000000000003F0F7FC30DC3F7FC00F7FDF0C3003ECDFDFC3DF5C3FF;
defparam sp_inst_3.INIT_RAM_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //t20k_romram
