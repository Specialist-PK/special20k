//Copyright (C)2014-2025 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.11.01 Education (64-bit)
//Part Number: GW2AR-LV18QN88C8/I7
//Device: GW2AR-18
//Device Version: C
//Created Time: Tue May  6 16:30:57 2025

module t20k_romram (dout, clk, oce, ce, reset, wre, ad, din);

output [7:0] dout;
input clk;
input oce;
input ce;
input reset;
input wre;
input [12:0] ad;
input [7:0] din;

wire [29:0] sp_inst_0_dout_w;
wire [29:0] sp_inst_1_dout_w;
wire [29:0] sp_inst_2_dout_w;
wire [29:0] sp_inst_3_dout_w;
wire gw_gnd;

assign gw_gnd = 1'b0;

SP sp_inst_0 (
    .DO({sp_inst_0_dout_w[29:0],dout[1:0]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[1:0]})
);

defparam sp_inst_0.READ_MODE = 1'b0;
defparam sp_inst_0.WRITE_MODE = 2'b00;
defparam sp_inst_0.BIT_WIDTH = 2;
defparam sp_inst_0.BLK_SEL = 3'b000;
defparam sp_inst_0.RESET_MODE = "SYNC";
defparam sp_inst_0.INIT_RAM_00 = 256'hE552E0B2CBC8D6F83577E2D9F6E2A8C82655557A2935555C7A07A41500FEAF4F;
defparam sp_inst_0.INIT_RAM_01 = 256'h9A27A9E6589E2499EA78B21F2041252C2CBA09959B4EFAD55095DDCDD9C88A74;
defparam sp_inst_0.INIT_RAM_02 = 256'hA77EED9518E7B6CBC8104017E96657E966597F96A1727C957E966497F9EA177B;
defparam sp_inst_0.INIT_RAM_03 = 256'hD7CB2696F9AADA15E6E2E9EECA9BAB685AF2B795FE551D89BD4595495546977E;
defparam sp_inst_0.INIT_RAM_04 = 256'hE5169BBB687B62F97E67EA5D1C958B4BFDBB1860A5EF65EA66EEDA1E6A4EEE3E;
defparam sp_inst_0.INIT_RAM_05 = 256'hBE7EF246FB2E991E8A157AE1B5BD0FC955564FA55CBF287B2FC8FBD5647D5D96;
defparam sp_inst_0.INIT_RAM_06 = 256'hB6C940004A225209FC13A3CBE5F94789561563763EBDF8A3476ACB22CBE172AC;
defparam sp_inst_0.INIT_RAM_07 = 256'hBF780157A41F9B07FA9BE2D54FF957EE96FBBA6CFEFAA7AEDB6D77ED8A2DBF9D;
defparam sp_inst_0.INIT_RAM_08 = 256'h0020021DB7EF8EA09BD7ED4117D04D0F342E4637E9D20BE42CDFD2FD2FD2FBF4;
defparam sp_inst_0.INIT_RAM_09 = 256'h00CEE4E40044E4E70089F9DE0088387600F0817900600D91316F83000CFA0C1A;
defparam sp_inst_0.INIT_RAM_0A = 256'h0024000000C0000000C0019002A02002002A19283C24098C2BBA002A00000000;
defparam sp_inst_0.INIT_RAM_0B = 256'h00960260033020020000000009D625960027258325632BAA25A7309620002576;
defparam sp_inst_0.INIT_RAM_0C = 256'h25561755155D340018092555200215D537060083308325562406259617582376;
defparam sp_inst_0.INIT_RAM_0D = 256'hC00000062AAA0600200230A70025162525550295255500032586189619560096;
defparam sp_inst_0.INIT_RAM_0E = 256'h255615D5155D155718091575157516250007035C30831EAA1EAA258317582556;
defparam sp_inst_0.INIT_RAM_0F = 256'hFFFF15D51D5525D6355525961555258025961595009500032406009615D71557;
defparam sp_inst_0.INIT_RAM_10 = 256'hA9EE288E22B86259AE217D565E4B37EB7607D2CB0477D30638E79E3EF38FFFCB;
defparam sp_inst_0.INIT_RAM_11 = 256'h76441F9107644A5752E717E7E415FEFE50547E50BA38BB6E2A92E698AA188AE4;
defparam sp_inst_0.INIT_RAM_12 = 256'h9F6FB6F41F9765FBD9AF4B757114799579076EBED5B9AF779657655465117B90;
defparam sp_inst_0.INIT_RAM_13 = 256'h6971979071C5E5E6F4A9E6F7BECB9C75975F9AD8FA8B5F90556BFAAD2D145907;
defparam sp_inst_0.INIT_RAM_14 = 256'h72526F5971AC1CA5D41FA5E41EA5C7D88D1E85FBCBEBF4BF4B5BFEADE6B5C6AF;
defparam sp_inst_0.INIT_RAM_15 = 256'hAFC8DC6C6C7C4C55C6B9E79AFC6AEC6A716EC6B9EA2D4B9B6B1E71C65D7E4155;
defparam sp_inst_0.INIT_RAM_16 = 256'h656D9726CF8A2C55F361287A127C97A0CF61DF6C8DDBE6C8BD472712EAF1317E;
defparam sp_inst_0.INIT_RAM_17 = 256'hF7A65ED0F6171E9C1CB6F07A7D957E77ACE6E9BCB69435EB97A557F1F9147E57;
defparam sp_inst_0.INIT_RAM_18 = 256'h14559656512FC35F65965965814EA3FC368BC352F0D7D965604A659656DF7755;
defparam sp_inst_0.INIT_RAM_19 = 256'hF87647E47647CAC47F652B43658686E389D0BDA2055DF18D0C1E138D76050597;
defparam sp_inst_0.INIT_RAM_1A = 256'h520E1F499E226889EA78BDC51715227A2E89B92A889DFF555D58868172DBF876;
defparam sp_inst_0.INIT_RAM_1B = 256'h8BA26E9AA62519F7FF67D5753D3F55625AA9F659607DF5574E1287A12D236749;
defparam sp_inst_0.INIT_RAM_1C = 256'hFB8B8BAABB2A5561652CEF4E86FF658B43659620584A7E10BA7975498749E61D;
defparam sp_inst_0.INIT_RAM_1D = 256'hB6EABAA53642C9656529798890E54BA6AE787E1FFD5878695639BBB685B93BB9;
defparam sp_inst_0.INIT_RAM_1E = 256'h8000011157160E2F0CB1B4A179F18696165A29572076727F2EBE7FBF88890552;
defparam sp_inst_0.INIT_RAM_1F = 256'h04C7050121041441C618500024FC6079F9136109A6F84D849819A089A0C49854;
defparam sp_inst_0.INIT_RAM_20 = 256'h34245E7B6ECFF0BE388EE3FC2A2BA97BA541645A05106519CA929421F2C51049;
defparam sp_inst_0.INIT_RAM_21 = 256'hA2BB43A54AE6D16C5BA4B06518A1481E14812189934EE351B9A42CA2B84998BF;
defparam sp_inst_0.INIT_RAM_22 = 256'h5A5585E76A9B439455CD6AAA6A188296D6B268A8461610E90DA4394E70D1B5AC;
defparam sp_inst_0.INIT_RAM_23 = 256'h7F18AA29BA62369AC5151445245451FE3EEEE45690534105EAB7BADE6B76A918;
defparam sp_inst_0.INIT_RAM_24 = 256'hE99A6A98A220AA2E2058AD2AB62A81D6279E288AA76F5996E5F148521496A571;
defparam sp_inst_0.INIT_RAM_25 = 256'h10508215402E4628F85163624030CC90E4FA21A47C7118E264941A5E36655FA6;
defparam sp_inst_0.INIT_RAM_26 = 256'hA5D079766B58AB5B66A4991AD297A612A56C931EE9841A5BEE2696929E9A9584;
defparam sp_inst_0.INIT_RAM_27 = 256'hA3268C9637A4A1AB907169A697A4A1A69A50757A2A6DAE9B560412ADEDAA9A69;
defparam sp_inst_0.INIT_RAM_28 = 256'h184669EA78A9A62D4A205618467E9FA48A75D62D5A205493D5F2462A85D4D527;
defparam sp_inst_0.INIT_RAM_29 = 256'h0004C3055353539C524D7CF7EFDCBDBEBF9CBDBEBF9BBB9F22624DD286E2B996;
defparam sp_inst_0.INIT_RAM_2A = 256'hF26B9AA5A92D9E78E1A5FCF9FCF19793F296969FE1AD05C356EEE6BCAF19FFF4;
defparam sp_inst_0.INIT_RAM_2B = 256'h952D17BE11B6AB6BA17967C8B5B9B6AA759D29A4BA56A23676F4F2D26896E569;
defparam sp_inst_0.INIT_RAM_2C = 256'h9BA258D861AB37776258D851B9526B68D85168194C919E2EA2919C13D418A541;
defparam sp_inst_0.INIT_RAM_2D = 256'h2CBCBCBDA5255961762665DB896E9BF66EA2EEE514A6A913613697481AA9429A;
defparam sp_inst_0.INIT_RAM_2E = 256'h566E2D5969EEA565869CB595C5559BD882F31C7EE62E12E1507EEE96262A4196;
defparam sp_inst_0.INIT_RAM_2F = 256'hBBE4537BE9F547FF64D767957EF22FAE4ED6F8A6E45B907B1515E9A3DC9EC91C;
defparam sp_inst_0.INIT_RAM_30 = 256'hE850A854799654B94A6424B9118B37BE5F4E6E05FB95723882D2388ACAAB2AAF;
defparam sp_inst_0.INIT_RAM_31 = 256'h000000000000F51E56E0539E56E84EA1464B911E6D179AE1D4715B81465C66C6;
defparam sp_inst_0.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_38 = 256'h86DE5E2982E26964E7DD265205EB499D264A6789665A2D9D6149295E6A2C1741;
defparam sp_inst_0.INIT_RAM_39 = 256'hE3DEEE629971C941E3DEEE66855B6AEEE1B88E7EB9A589AE882E5E6BA60B0BB9;
defparam sp_inst_0.INIT_RAM_3A = 256'hDA6899758F169DA4B95E66B5A89B7B895296EB89EE52DE7E9979AEEE69B9791E;
defparam sp_inst_0.INIT_RAM_3B = 256'h0035A2094D16A92685616B9A64B053E8F23C8F62E10512E5BBBBE9A299EE2169;
defparam sp_inst_0.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_0.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_1 (
    .DO({sp_inst_1_dout_w[29:0],dout[3:2]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[3:2]})
);

defparam sp_inst_1.READ_MODE = 1'b0;
defparam sp_inst_1.WRITE_MODE = 2'b00;
defparam sp_inst_1.BIT_WIDTH = 2;
defparam sp_inst_1.BLK_SEL = 3'b000;
defparam sp_inst_1.RESET_MODE = "SYNC";
defparam sp_inst_1.INIT_RAM_00 = 256'h8EA1E27847F7C7C72AB761E2BC103FF8639560B600A555503A03480505303F00;
defparam sp_inst_1.INIT_RAM_01 = 256'hCAF1ACAB3AC6B2BC2B18FE03C2030F231F3911F8E78C7AE0031D439438EA4444;
defparam sp_inst_1.INIT_RAM_02 = 256'hB3F0BC952C2BFACCF080C00CE4C7CCE4E3F4C44A3CC1103CCE407C4C440FCC1B;
defparam sp_inst_1.INIT_RAM_03 = 256'hC4D3E2123401C87104F1C8CFC8B28721C2760F540F603C0D100D5A01600113F0;
defparam sp_inst_1.INIT_RAM_04 = 256'h8C3523C721FC23F9B03B03103D20D745561BFC811E5F210044F1C87D8ABBF48D;
defparam sp_inst_1.INIT_RAM_05 = 256'h86BE7663F3020C338C30F8C30C7802FA55801FA58F2BE3FFC0F9B78603786FA0;
defparam sp_inst_1.INIT_RAM_06 = 256'h724D40008C83218C2002C0CBC8030F4E00B5482C8E3C13C80C2BD3C1F80202BF;
defparam sp_inst_1.INIT_RAM_07 = 256'hF1FC02004DBC0E6FC3456B5501FA0B2019C3C0B330C078C6C722F0685A3CB76C;
defparam sp_inst_1.INIT_RAM_08 = 256'h020800EC88FF1EB8BC7B22DB7FC510601E3F9C5C0EB2D4F941747B47BC7BC11E;
defparam sp_inst_1.INIT_RAM_09 = 256'h00FA550000CA550200AB9D9200F5F01900FC26CC00E88AAC330703E0033E0C06;
defparam sp_inst_1.INIT_RAM_0A = 256'h02403C0000C027C005D405D4240606A4004531E9024A1DDD2BBA002A11550000;
defparam sp_inst_1.INIT_RAM_0B = 256'h110324060330062427CF3C3C30C330C32A4330C93033032430433243355D3243;
defparam sp_inst_1.INIT_RAM_0C = 256'h300300600058300001903000355700C0300300C330C33AAB300330C303093143;
defparam sp_inst_1.INIT_RAM_0D = 256'hC0000003300300603AAB32C315600260254016803000155730C301C3310300C3;
defparam sp_inst_1.INIT_RAM_0E = 256'h300300C000582AA901900241024002600003175D30C30EA90C0030C3030905D4;
defparam sp_inst_1.INIT_RAM_0F = 256'hFFFF00C00D55304335543043258030C030C305D409801557300300C309C30003;
defparam sp_inst_1.INIT_RAM_10 = 256'h8EA79AFA7EAFEFDBFE7CF3EFFC24AF8F3083C82C0B8A200ACF3CF3CA00E04124;
defparam sp_inst_1.INIT_RAM_11 = 256'hF6AFFDABFFEAECC8D7D34BAB8BF81EFBBFE6C378FF48BE23C9E678AF6FAAF638;
defparam sp_inst_1.INIT_RAM_12 = 256'h87ADB4080C0701F2F230A49C22BAC6BB38238DF4989AC6A0FFB6BF8AFFAB6E6F;
defparam sp_inst_1.INIT_RAM_13 = 256'h2FF0FFC5F0C28E8B1ECE8B1FF0C6BC30FF0F2A7A3CA98C23B568F2A792BAEB23;
defparam sp_inst_1.INIT_RAM_14 = 256'hBE8DDC1FFC83FFBFE3FCBFD3FEBFC33B172EBBCAF2E11EF1ECBA02A68AF0C2A7;
defparam sp_inst_1.INIT_RAM_15 = 256'h808970F0E0E0F0F00DEFBEF900E27C28C3B30DEFF22606B0FF0AF0C3FC308ED5;
defparam sp_inst_1.INIT_RAM_16 = 256'hA03E2E8F3B3F3C166C3BBEFFBB6BAE8BB03BD76B97D2EF8AC7DA0C33F803C3F2;
defparam sp_inst_1.INIT_RAM_17 = 256'hCE4F7FF07ABF4B13F57AAFECEE956043C34BF9DC3AFE5CF38788003CE3EDF656;
defparam sp_inst_1.INIT_RAM_18 = 256'h07B8EFFFFDD025CCFFFE4EFFFF72EE025CF025CD09733FFF7FFAB8EFF7B02C00;
defparam sp_inst_1.INIT_RAM_19 = 256'hD0B4CF0CF0CCC2C3CCFFC065FBEFFAFD8ECF9DB1FE220E17F3378E977302FCFF;
defparam sp_inst_1.INIT_RAM_1A = 256'hF4B3BDCBF6BFE3C70BC8C7C17706119747D8F76BD8E3036ABBEBEF80B2CAC9F6;
defparam sp_inst_1.INIT_RAM_1B = 256'hD1F63DEAFA383B1D55EC77878B81CFEBEAF71FBFFFF3EE01D3BBEFFBBB65F8D2;
defparam sp_inst_1.INIT_RAM_1C = 256'h3D2BC72C3F22D6077790F1CFFFCCFFD065FBFF1FEECFC3B8FF8FF884EF4653BD;
defparam sp_inst_1.INIT_RAM_1D = 256'hFECAF2BA1F1BFA3737BDFDC8C3798576BDBFE7FFFE0EEEEFD4813C721EDAEF7D;
defparam sp_inst_1.INIT_RAM_1E = 256'hC0000330F403BC7E0C36FCA022B2EEE3BB6B2E03C23C70C13EBCC181AC48015B;
defparam sp_inst_1.INIT_RAM_1F = 256'h0C0C0EEB23CE34D30C34C00035D48022BB30440AF7E8C110AECCE0B860C38438;
defparam sp_inst_1.INIT_RAM_20 = 256'h4846B3A0D30C001328CA61000E19F819C0480EBFAF0ACC33078B7CC281420ACC;
defparam sp_inst_1.INIT_RAM_21 = 256'hA3CE2800807C39FA7F1C4AC0287ACC71ACC79224E200FAD09310C4E38F0BEE73;
defparam sp_inst_1.INIT_RAM_22 = 256'h3E132085FF80E832F02338EE327DAA00300F38FF028FC003000E8304EA300CC4;
defparam sp_inst_1.INIT_RAM_23 = 256'hF1BC4EB1BC6B8F802F9E9E2BF67E7D86B13132F7810C40008FC23F08FC5FF80A;
defparam sp_inst_1.INIT_RAM_24 = 256'h708C6B08423BC232102D0BB02F4C00A00C00330EB4301BC6712AEEB3AEC6BC4A;
defparam sp_inst_1.INIT_RAM_25 = 256'h002080B8800F80F13C22111002110824FC232304EC89E4F22CBAB224082AAD40;
defparam sp_inst_1.INIT_RAM_26 = 256'h0E4ACC4232CCD2CCE33EC80CB33C04B10E131E28C3C002DC27B0BCBCB8B8B62C;
defparam sp_inst_1.INIT_RAM_27 = 256'h142C50B1493CC0C3CACC430C393CC00C30CAC44C10CBB38C3B00034B702C30C3;
defparam sp_inst_1.INIT_RAM_28 = 256'hB2DC4B32CC4BF020EC25D8B2D044310C4F0BC020CC25D8DDEAD19E3CA02CC52E;
defparam sp_inst_1.INIT_RAM_29 = 256'h3139041786C6D61D37DB9EF9EDA6CEC6CCE6C6C6C4E4C4E01CE6D7E7C331CE48;
defparam sp_inst_1.INIT_RAM_2A = 256'h037BDEB5BD65BBB4B8E40259425AE60A01A7173065E6126F391139A86A1F0009;
defparam sp_inst_1.INIT_RAM_2B = 256'h515200034AC72C72F4998C0CE419C5BE94312DA4D190F196C507231469DABA53;
defparam sp_inst_1.INIT_RAM_2C = 256'hC0F0B93E34F1FBBBBC893D2C63A2BA993C2CBAB60539FEAA61B9F8013C44922B;
defparam sp_inst_1.INIT_RAM_2D = 256'h26CEC6CCFC017E389105FC71E9BCF1FBC92C593A087E49F6F04FCBC0CC147DEA;
defparam sp_inst_1.INIT_RAM_2E = 256'hD34F8D7F3453E5F8D1371C9A82AAD358F1F938187651F51F84EB13E38F25DBE3;
defparam sp_inst_1.INIT_RAM_2F = 256'h1D3C0000344D6355388561352090D1E6663073693844E11C817579F94631CD87;
defparam sp_inst_1.INIT_RAM_30 = 256'h00180E46EC97CDC9207E67C98AE30003C4E4F0027184CD9BEA30B3C7A8F8B3E6;
defparam sp_inst_1.INIT_RAM_31 = 256'h0000000000020585D3002805D300243A227C98AB09B2CB0B16134C00AC04F083;
defparam sp_inst_1.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_38 = 256'hB67EC34EBA72C2DF04C7EDFE034BFB77EDFC3F9F2DF61CBF7AFFCD3CF30EBE00;
defparam sp_inst_1.INIT_RAM_39 = 256'h6F336B6DC2BCC7846F336B6F35C1FB093D1CBC40ECB8C0F0EB8FC32C3AE13D9C;
defparam sp_inst_1.INIT_RAM_3A = 256'hF7C1F7FDF0AEFF7F2E3C3F2FCBCAE1C83CE30EC3CB3CBC40DE2DB093B8D9DBB4;
defparam sp_inst_1.INIT_RAM_3B = 256'h0021030B5FAC84200028E0B810A01E3F87E0F8792FAF492BCADB0DB4EB272AFF;
defparam sp_inst_1.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_1.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_2 (
    .DO({sp_inst_2_dout_w[29:0],dout[5:4]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[5:4]})
);

defparam sp_inst_2.READ_MODE = 1'b0;
defparam sp_inst_2.WRITE_MODE = 2'b00;
defparam sp_inst_2.BIT_WIDTH = 2;
defparam sp_inst_2.BLK_SEL = 3'b000;
defparam sp_inst_2.RESET_MODE = "SYNC";
defparam sp_inst_2.INIT_RAM_00 = 256'hCEB2900E903B130B2AA0A92F8F037F385BF188CE23CAAAA00E0CEC2200333FC0;
defparam sp_inst_2.INIT_RAM_01 = 256'hC4301CC720C0720C4302CE00E084080323E007F3CAC8CF09300AC8EC8D380C18;
defparam sp_inst_2.INIT_RAM_02 = 256'h303333A3088FCB0438210004805FC48457F8484D3C4210204809FC84805FC411;
defparam sp_inst_2.INIT_RAM_03 = 256'h8C3CB00030C2CC4300FFCCCFCC400B3108CF03088788C3CE001100100C832033;
defparam sp_inst_2.INIT_RAM_04 = 256'h804423CF3130032C33733330C3C8CAE00334300820EB33040CF3CC4C818CE80E;
defparam sp_inst_2.INIT_RAM_05 = 256'hC886CFDB2CF04CC00CC30B8800CA123BC62C50BE03A8E310EA3BBCA084CAA280;
defparam sp_inst_2.INIT_RAM_06 = 256'hB34100001813C94F2020CC3CB00013101809002003BE10C020CF3CB02C80C8F2;
defparam sp_inst_2.INIT_RAM_07 = 256'hE33C001C400CCB01CCC93074103C18F0113FC0730F8CBCFF4B300C0C853CC3B4;
defparam sp_inst_2.INIT_RAM_08 = 256'h018000E28CF3C8300CC8A30C20414E32303308208CF3C4F0488CC34C34C32A30;
defparam sp_inst_2.INIT_RAM_09 = 256'h0040000000BFFFFF00EFEABA00BEAFBE00EABEBF00042450381059E0000F2687;
defparam sp_inst_2.INIT_RAM_0A = 256'h0400000000400000004001100000000000000500040504100110000000000000;
defparam sp_inst_2.INIT_RAM_0B = 256'h0004000001100040000000001014051400010550041501400401140400000554;
defparam sp_inst_2.INIT_RAM_0C = 256'h0554155515551555155505000000155505541555155510010554155515500554;
defparam sp_inst_2.INIT_RAM_0D = 256'h4000000400000004000014010005140505550015055500010414155505541555;
defparam sp_inst_2.INIT_RAM_0E = 256'h0554155515551000155515551555140515550154155514000555155515501555;
defparam sp_inst_2.INIT_RAM_0F = 256'hFFFF005505550404155504041555155515551515101500010554155510141555;
defparam sp_inst_2.INIT_RAM_10 = 256'h1C4711CC730C8320C8320000418C00AF8A0BF10000010400C10410410400C30C;
defparam sp_inst_2.INIT_RAM_11 = 256'h0A108184206104000014A0A0A0865B6C82188880CC400C8730C8330C4330C031;
defparam sp_inst_2.INIT_RAM_12 = 256'h6C718AAC22ACA81A18768C12EC410C4105387FC6A13C8F22108204C104C42202;
defparam sp_inst_2.INIT_RAM_13 = 256'h310E10210138400730C00733CF8C41421023CCF10F13C1A801843C4F30410434;
defparam sp_inst_2.INIT_RAM_14 = 256'h0E233CA10E30808428828418808428020850802A0A0A30E30CC0184C0D01384C;
defparam sp_inst_2.INIT_RAM_15 = 256'h320081313131313912C000002104F38C047012C03CCF0E123CE101384086A006;
defparam sp_inst_2.INIT_RAM_16 = 256'h4830F083822F0288C400003000213C0F12000C71081C4300CC004043C304C4C6;
defparam sp_inst_2.INIT_RAM_17 = 256'h00C484700320E1080003A200E0F18C28280F0A01C3002208283E4EC20F200218;
defparam sp_inst_2.INIT_RAM_18 = 256'hA000204C4C00820000100204C808C30820CC8231208000043208F02043128493;
defparam sp_inst_2.INIT_RAM_19 = 256'h0A82102102100C2080003202080201F06F2330C420C8F2080080F208C3002210;
defparam sp_inst_2.INIT_RAM_1A = 256'hC4F80320C03B23D09B26CC0054A8D7345314D81F16C0422A8822C302030A0802;
defparam sp_inst_2.INIT_RAM_1B = 256'h14C53607C5B0C8300020C040888B100301C43081320030931000030008420413;
defparam sp_inst_2.INIT_RAM_1C = 256'h3A03FF303F3108C4C8307307108000320208134200204800CC41023700DCDC03;
defparam sp_inst_2.INIT_RAM_1D = 256'hCF01C03C30DF3CC808023026CC3F3001321334C00440000204033CF3120633A0;
defparam sp_inst_2.INIT_RAM_1E = 256'hAAAAA83AAFBAEBEA2EEEAA82AAE8000004040F90E380081B43C01B5B73114867;
defparam sp_inst_2.INIT_RAM_1F = 256'h0D4C4E08830C30C30C30C2AAAABEBEAAE03BBAABBAA0EEEABBAE82EA82EAAAE8;
defparam sp_inst_2.INIT_RAM_20 = 256'h11C008A5199CA63B62D8D4258D53D963D296600C112116508DAC410F2301211E;
defparam sp_inst_2.INIT_RAM_21 = 256'hCBE6846A197141384E4D811251B021C0021C060AC018F12754754D0B56403B54;
defparam sp_inst_2.INIT_RAM_22 = 256'hC65475D421A50469061C51D652048579072B70F69D719018426047972112510D;
defparam sp_inst_2.INIT_RAM_23 = 256'h0B0CD4741D0301A610131300804C4E81C4B99909A014A00983E60F983E421A75;
defparam sp_inst_2.INIT_RAM_24 = 256'h75DD335F58B2D4350084945251248285C141B70D057260D8F62000080018BD80;
defparam sp_inst_2.INIT_RAM_25 = 256'h108CC182033F33360C5061616170104200462050009802030000458D815AA057;
defparam sp_inst_2.INIT_RAM_26 = 256'h70F11AD83700E701C3700A0DC051018460163E7D1C28161D833D8D8D8D8D8F60;
defparam sp_inst_2.INIT_RAM_27 = 256'hD103440D1371026FE11E9C71C3710271C7211E90271CC40D0804239CC62DC71C;
defparam sp_inst_2.INIT_RAM_28 = 256'h861818B62C18F9D411D42186102DCB700F98C5D411D420A52CF15436D860D102;
defparam sp_inst_2.INIT_RAM_29 = 256'h01138E1C342626718514030D34C0E0E4E4CCECECECC2264429051487C3B0EDE1;
defparam sp_inst_2.INIT_RAM_2A = 256'h9373D4B42D4D4019F6D524F508F3C73C91460609D18F009E73BBB1645910A950;
defparam sp_inst_2.INIT_RAM_2B = 256'h4B612EED63E63E63D635024ED535C62D37090D42C1DCB43516171B5454D03C60;
defparam sp_inst_2.INIT_RAM_2C = 256'h5CD74D44504A88889259445443574A59445448448D0581392585801370403CC4;
defparam sp_inst_2.INIT_RAM_2D = 256'h71E1E5E5D6018591398516435E165AA1690E3D951896454712616248659673DF;
defparam sp_inst_2.INIT_RAM_2E = 256'h15B9798599713616450634D146AA6E45F2A5849CDB510610272899597D751459;
defparam sp_inst_2.INIT_RAM_2F = 256'h3CB49EEEDA605700B41991466550550D4D5371519412115C198972F3E40BA256;
defparam sp_inst_2.INIT_RAM_30 = 256'hA0854F8626A520685951CF6A3C5EEEED66151A0873552761F61341CF98B552D7;
defparam sp_inst_2.INIT_RAM_31 = 256'h000000000001C04609A0874609A0953C90F6A3C9A98A69A40118268211861A49;
defparam sp_inst_2.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_38 = 256'hD0DF4134DCD37341420DC41E01CE7105C414360D04182CD47031E49F7D3846A3;
defparam sp_inst_2.INIT_RAM_39 = 256'hDE79292C493C8B009E792927F1437D299434D819E4914CD34D8F4124925074C4;
defparam sp_inst_2.INIT_RAM_3A = 256'h4370D051D8021437A45F353D4F4A534D1E493E4DCFDE9419C4A49299514857D4;
defparam sp_inst_2.INIT_RAM_3B = 256'h00004B2C00460A38C63143D428D05521445114030811E3084A48A4934D4D3031;
defparam sp_inst_2.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_2.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

SP sp_inst_3 (
    .DO({sp_inst_3_dout_w[29:0],dout[7:6]}),
    .CLK(clk),
    .OCE(oce),
    .CE(ce),
    .RESET(reset),
    .WRE(wre),
    .BLKSEL({gw_gnd,gw_gnd,gw_gnd}),
    .AD({ad[12:0],gw_gnd}),
    .DI({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,din[7:6]})
);

defparam sp_inst_3.READ_MODE = 1'b0;
defparam sp_inst_3.WRITE_MODE = 2'b00;
defparam sp_inst_3.BIT_WIDTH = 2;
defparam sp_inst_3.BLK_SEL = 3'b000;
defparam sp_inst_3.RESET_MODE = "SYNC";
defparam sp_inst_3.INIT_RAM_00 = 256'h7010402C6C3D604D301AC3B1EC3EEDB3F37FFFECCE4FFFF02CC2C00F0DF08733;
defparam sp_inst_3.INIT_RAM_01 = 256'hF73DCF33CCF33CCF33CCECDEC03333DD0B13FFDE787BAC7FFEC0774777B0370F;
defparam sp_inst_3.INIT_RAM_02 = 256'h0EF00B3F3BB5EC7BB00CC0374F7F774F736374F33770DCCF74F3F4374F3B77DC;
defparam sp_inst_3.INIT_RAM_03 = 256'h7BB2CFCFF3F3C37EF3FFC3FFC37DCF0DFFACEF3FB4FF7B13EFEC3FEC7FCDCEF0;
defparam sp_inst_3.INIT_RAM_04 = 256'h73B0DFCF0DF37BB3F08F08EF7B3F71AC01CC30F7CFF30EF333F3C37C730CC73C;
defparam sp_inst_3.INIT_RAM_05 = 256'h37ECACF3B2CCEF7DEFBEECB7EC2CDFB1FFFFB2CFFB02CED2C0B032CFFB2CFB3F;
defparam sp_inst_3.INIT_RAM_06 = 256'hF043C000CFF7F3DFCC0EFFB2CFDCEF03FFFFFFEFFB3CDEFFEF33B2CBB333F73B;
defparam sp_inst_3.INIT_RAM_07 = 256'h1DF003FFF3BC0DEDC0CD107FEDB3FACEC0B33B3EECBBF7B94F0FDBB8F7BC11D4;
defparam sp_inst_3.INIT_RAM_08 = 256'h00BF33FB37CB373CCF3ECFF3CECE34CCCF35F3CC079E73CF333770770770B1DC;
defparam sp_inst_3.INIT_RAM_09 = 256'h002A00000000000000155555001555550041555500020002015550000FEC0438;
defparam sp_inst_3.INIT_RAM_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_10 = 256'hDFB7FDF37DDFB7EDF37FF7DF3D33DE872CC1CFFF0FBEFB0F7DF3EF7CFFFF7CF3;
defparam sp_inst_3.INIT_RAM_11 = 256'hE8CF7A33DE8CFF3CF0F28E8E8F7311473DCFB3FCD73EDF77CDF37EDF37EDF77E;
defparam sp_inst_3.INIT_RAM_12 = 256'h868A28000A3E8FA3A310F3DF477DF37D28028C68FDE739FCCF3FFB7CFB73C47D;
defparam sp_inst_3.INIT_RAM_13 = 256'hCCE8CF8CECA3F3FFDC03FFDF2C833B2CCF8B3B9FECFE7A17BFF3B339CF7DF702;
defparam sp_inst_3.INIT_RAM_14 = 256'hECF00C3CF8DF7A33E37B33E37A33D37DF35A3BB3A3A1DC1DC3FCC33BF86CA33A;
defparam sp_inst_3.INIT_RAM_15 = 256'hFCCF3FDFDFDFDFDFFF33CF3FCFFF9A3B3FC0FF33B3B9C0EC368CECA33E285EFF;
defparam sp_inst_3.INIT_RAM_16 = 256'hBF3A13730DCD093F73FF0FD3F0CCE779CCFF768CF3A373DCF35F33F0CDFF7F68;
defparam sp_inst_3.INIT_RAM_17 = 256'hDFF3F44A68EF4FC334E80DFF0A3FFB0E8339A35A28DFCFA28E87F468A1FD68FF;
defparam sp_inst_3.INIT_RAM_18 = 256'h4FBFCFB7B7DC3CFDF7ECFCFB77F78CC3CC733CDCCF3F7DFBDDF39FCFBDECFBFF;
defparam sp_inst_3.INIT_RAM_19 = 256'hA168CE8CE8CCA093BDF7EC3CF3FC3F7FCD6EEA10DFF30EF3EFB67EF3D903DFCF;
defparam sp_inst_3.INIT_RAM_1A = 256'h7793F5ECFB30DCCF73DCF3A35E4F33CF37CDDF73CCF3318033CCF300E8A3A168;
defparam sp_inst_3.INIT_RAM_1B = 256'hCDF377CCF73FBFCD00FF3FFFB3B1FFF3FCF7CF3EDDF7CFFDDFF0FD3F037CF7DE;
defparam sp_inst_3.INIT_RAM_1C = 256'hF1DFFF0EFF0DFFF7F7CF3CF3DF3DF7CC3CF3ED0DFFC333FCD77CF4CFFDCF3FF7;
defparam sp_inst_3.INIT_RAM_1D = 256'hECCCF337CFFFB3FFFF0FD3FCF737CCFF33DED7B007FFDFDEFF7CFCF0DDEC331E;
defparam sp_inst_3.INIT_RAM_1E = 256'h0000000155155555005554005553FC3FF0F0CDFEC33333010B330101102083FE;
defparam sp_inst_3.INIT_RAM_1F = 256'h0141405100410410410410000554545550015505555005545555401540055454;
defparam sp_inst_3.INIT_RAM_20 = 256'h5F7331FED1330DE1DCF78DC378DE70DE7CF0FF30CF0CF8CC0300CF3900030CF4;
defparam sp_inst_3.INIT_RAM_21 = 256'hF34C33E3FBDFBCD33537FCFCFCDCC370CC370FCF403BFCFFF7E3BBB30C004055;
defparam sp_inst_3.INIT_RAM_22 = 256'h3C37E37DC30EF3E37DFBDDCC345D33E37CC3CCDC3FCF0CFFCFFF3E3EFCF0EF3B;
defparam sp_inst_3.INIT_RAM_23 = 256'hD1CC333CDF33CF0FF7CDCDF30F3737C659111F7F003FC0C3B74EDD3B74DC30FF;
defparam sp_inst_3.INIT_RAM_24 = 256'h3ECFB3ECF73CFB30003D37F4DF4D00FF30DC0CCC0CFCFCFF9FCCC330CC3F37FC;
defparam sp_inst_3.INIT_RAM_25 = 256'h003C03FFC30CF00FC0C1C1C1C1F178545054005414115450400F3E3373B004FB;
defparam sp_inst_3.INIT_RAM_26 = 256'hFFBCFCF73FD3FFD373FD08CFF4FF73F0FF3CE4DA7F428FE3387FF7F7F7F7FDFC;
defparam sp_inst_3.INIT_RAM_27 = 256'h150054015EFD00D33CFCFFFFFEFD00FFFFFCFCFF7FFF4ECF34400FFF4DEFFFFF;
defparam sp_inst_3.INIT_RAM_28 = 256'hFFF73F1FC43FCFFCD3FCFFFFF707F1FC3FF3C3FCD3FCFC158700733D3FCCCF00;
defparam sp_inst_3.INIT_RAM_29 = 256'hCCCC30FFFFFEFFF3FFFFD965967646464676464646744470048EFBB7771DC70F;
defparam sp_inst_3.INIT_RAM_2A = 256'h0EDCFB3ECFBB70FF7DCDC393732E7CE40E3CCCC0433903659E221E0380F3000C;
defparam sp_inst_3.INIT_RAM_2B = 256'hC3CF04470E4FE4FE70E3F0380FE37DCCEEC3FBB0137B30EDCDCDC03BECFF37DC;
defparam sp_inst_3.INIT_RAM_2C = 256'hC330C3BC30C1622230C3BC30DC30C3C3BC30C33C33BFF7CFCF3FF40CCC5403F3;
defparam sp_inst_3.INIT_RAM_2D = 256'h0646464670033C30CFFCF0CEC3F0C16F0FF235130030FFFEF0EF0EC04C38FCF0;
defparam sp_inst_3.INIT_RAM_2E = 256'hFF0B0B3C30DF0CF0C3FDEC3CC000C2DCC06F3C33B0DFFCFFFFC111C3030EFFC3;
defparam sp_inst_3.INIT_RAM_2F = 256'hE51C344470EFFC00D00FFF7FF03F73F8F830EDCD10044037FF7FDFDCBEC283FC;
defparam sp_inst_3.INIT_RAM_30 = 256'h003ECDFCFC3CF5C3FBCF79C3E7C244470EFDF003EE3DC4CDDCF0CDC13330CCCF;
defparam sp_inst_3.INIT_RAM_31 = 256'h000000000003B0FCFF003EFCFF003F37FF9C3E7F0F3FC30DC3F3FC00F7FCF0C3;
defparam sp_inst_3.INIT_RAM_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_38 = 256'h3FBCDF0C37B0EEFF7067BFFC83B8EFF7BFF33DCFFFFBBC3F0CC3CC3CF30B3F30;
defparam sp_inst_3.INIT_RAM_39 = 256'hA5930F04C03C6D0065930F0F0FDEF30D1FEC3B007C30C030E3B7DF0C30ED8C1C;
defparam sp_inst_3.INIT_RAM_3A = 256'hF0ECFFFC33CC3F0F3C3C0DE779C3DEC3FCC307C337FCF3007C3C30D130C1CE73;
defparam sp_inst_3.INIT_RAM_3B = 256'h00155001557FCF0C3F0FFE7F3C083CC334CD334CF7CFCCF3C3C2CC30C3BB0CC3;
defparam sp_inst_3.INIT_RAM_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam sp_inst_3.INIT_RAM_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

endmodule //t20k_romram
